*Fully-connected Classifier
.lib './models' ptm14hp
.include diff1.sp
.include diff2.sp
.include diff3.sp
.include 'neuron.sp'
.option ingold=2 artist=2 psf=2
.OPTION DELMAX=1NS
.option probe
.probe v(output0) 
.op
.PARAM VddVal=0.800000
.PARAM VssVal=-0.800000
.PARAM tsampling=4.000000n
.include 'layer1.sp'
.include 'layer2.sp'
.include 'layer3.sp'
Xlayer1 vdd vss 0 in0 in1 in2 in3 in4 in5 in6 in7 in8 in9 in10 in11 in12 in13 in14 in15 in16 in17 in18 in19 in20 in21 in22 in23 in24 in25 in26 in27 in28 in29 in30 in31 in32 in33 in34 in35 in36 in37 in38 in39 in40 in41 in42 in43 in44 in45 in46 in47 in48 in49 in50 in51 in52 in53 in54 in55 in56 in57 in58 in59 in60 in61 in62 in63 in64 in65 in66 in67 in68 in69 in70 in71 in72 in73 in74 in75 in76 in77 in78 in79 in80 in81 in82 in83 in84 in85 in86 in87 in88 in89 in90 in91 in92 in93 in94 in95 in96 in97 in98 in99 in100 in101 in102 in103 in104 in105 in106 in107 in108 in109 in110 in111 in112 in113 in114 in115 in116 in117 in118 in119 in120 in121 in122 in123 in124 in125 in126 in127 in128 in129 in130 in131 in132 in133 in134 in135 in136 in137 in138 in139 in140 in141 in142 in143 in144 in145 in146 in147 in148 in149 in150 in151 in152 in153 in154 in155 in156 in157 in158 in159 in160 in161 in162 in163 in164 in165 in166 in167 in168 in169 in170 in171 in172 in173 in174 in175 in176 in177 in178 in179 in180 in181 in182 in183 in184 in185 in186 in187 in188 in189 in190 in191 in192 in193 in194 in195 in196 in197 in198 in199 in200 in201 in202 in203 in204 in205 in206 in207 in208 in209 in210 in211 in212 in213 in214 in215 in216 in217 in218 in219 in220 in221 in222 in223 in224 in225 in226 in227 in228 in229 in230 in231 in232 in233 in234 in235 in236 in237 in238 in239 in240 in241 in242 in243 in244 in245 in246 in247 in248 in249 in250 in251 in252 in253 in254 in255 in256 in257 in258 in259 in260 in261 in262 in263 in264 in265 in266 in267 in268 in269 in270 in271 in272 in273 in274 in275 in276 in277 in278 in279 in280 in281 in282 in283 in284 in285 in286 in287 in288 in289 in290 in291 in292 in293 in294 in295 in296 in297 in298 in299 in300 in301 in302 in303 in304 in305 in306 in307 in308 in309 in310 in311 in312 in313 in314 in315 in316 in317 in318 in319 in320 in321 in322 in323 in324 in325 in326 in327 in328 in329 in330 in331 in332 in333 in334 in335 in336 in337 in338 in339 in340 in341 in342 in343 in344 in345 in346 in347 in348 in349 in350 in351 in352 in353 in354 in355 in356 in357 in358 in359 in360 in361 in362 in363 in364 in365 in366 in367 in368 in369 in370 in371 in372 in373 in374 in375 in376 in377 in378 in379 in380 in381 in382 in383 in384 in385 in386 in387 in388 in389 in390 in391 in392 in393 in394 in395 in396 in397 in398 in399 out1_0 out1_1 out1_2 out1_3 out1_4 out1_5 out1_6 out1_7 out1_8 out1_9 out1_10 out1_11 out1_12 out1_13 out1_14 out1_15 out1_16 out1_17 out1_18 out1_19 out1_20 out1_21 out1_22 out1_23 out1_24 out1_25 out1_26 out1_27 out1_28 out1_29 out1_30 out1_31 out1_32 out1_33 out1_34 out1_35 out1_36 out1_37 out1_38 out1_39 out1_40 out1_41 out1_42 out1_43 out1_44 out1_45 out1_46 out1_47 out1_48 out1_49 out1_50 out1_51 out1_52 out1_53 out1_54 out1_55 out1_56 out1_57 out1_58 out1_59 out1_60 out1_61 out1_62 out1_63 out1_64 out1_65 out1_66 out1_67 out1_68 out1_69 out1_70 out1_71 out1_72 out1_73 out1_74 out1_75 out1_76 out1_77 out1_78 out1_79 out1_80 out1_81 out1_82 out1_83 out1_84 out1_85 out1_86 out1_87 out1_88 out1_89 out1_90 out1_91 out1_92 out1_93 out1_94 out1_95 out1_96 out1_97 out1_98 out1_99 out1_100 out1_101 out1_102 out1_103 out1_104 out1_105 out1_106 out1_107 out1_108 out1_109 out1_110 out1_111 out1_112 out1_113 out1_114 out1_115 out1_116 out1_117 out1_118 out1_119 layer1


Xlayer2 vdd vss 0 out1_0 out1_1 out1_2 out1_3 out1_4 out1_5 out1_6 out1_7 out1_8 out1_9 out1_10 out1_11 out1_12 out1_13 out1_14 out1_15 out1_16 out1_17 out1_18 out1_19 out1_20 out1_21 out1_22 out1_23 out1_24 out1_25 out1_26 out1_27 out1_28 out1_29 out1_30 out1_31 out1_32 out1_33 out1_34 out1_35 out1_36 out1_37 out1_38 out1_39 out1_40 out1_41 out1_42 out1_43 out1_44 out1_45 out1_46 out1_47 out1_48 out1_49 out1_50 out1_51 out1_52 out1_53 out1_54 out1_55 out1_56 out1_57 out1_58 out1_59 out1_60 out1_61 out1_62 out1_63 out1_64 out1_65 out1_66 out1_67 out1_68 out1_69 out1_70 out1_71 out1_72 out1_73 out1_74 out1_75 out1_76 out1_77 out1_78 out1_79 out1_80 out1_81 out1_82 out1_83 out1_84 out1_85 out1_86 out1_87 out1_88 out1_89 out1_90 out1_91 out1_92 out1_93 out1_94 out1_95 out1_96 out1_97 out1_98 out1_99 out1_100 out1_101 out1_102 out1_103 out1_104 out1_105 out1_106 out1_107 out1_108 out1_109 out1_110 out1_111 out1_112 out1_113 out1_114 out1_115 out1_116 out1_117 out1_118 out1_119 out2_0 out2_1 out2_2 out2_3 out2_4 out2_5 out2_6 out2_7 out2_8 out2_9 out2_10 out2_11 out2_12 out2_13 out2_14 out2_15 out2_16 out2_17 out2_18 out2_19 out2_20 out2_21 out2_22 out2_23 out2_24 out2_25 out2_26 out2_27 out2_28 out2_29 out2_30 out2_31 out2_32 out2_33 out2_34 out2_35 out2_36 out2_37 out2_38 out2_39 out2_40 out2_41 out2_42 out2_43 out2_44 out2_45 out2_46 out2_47 out2_48 out2_49 out2_50 out2_51 out2_52 out2_53 out2_54 out2_55 out2_56 out2_57 out2_58 out2_59 out2_60 out2_61 out2_62 out2_63 out2_64 out2_65 out2_66 out2_67 out2_68 out2_69 out2_70 out2_71 out2_72 out2_73 out2_74 out2_75 out2_76 out2_77 out2_78 out2_79 out2_80 out2_81 out2_82 out2_83 layer2


Xlayer3 vdd vss 0 out2_0 out2_1 out2_2 out2_3 out2_4 out2_5 out2_6 out2_7 out2_8 out2_9 out2_10 out2_11 out2_12 out2_13 out2_14 out2_15 out2_16 out2_17 out2_18 out2_19 out2_20 out2_21 out2_22 out2_23 out2_24 out2_25 out2_26 out2_27 out2_28 out2_29 out2_30 out2_31 out2_32 out2_33 out2_34 out2_35 out2_36 out2_37 out2_38 out2_39 out2_40 out2_41 out2_42 out2_43 out2_44 out2_45 out2_46 out2_47 out2_48 out2_49 out2_50 out2_51 out2_52 out2_53 out2_54 out2_55 out2_56 out2_57 out2_58 out2_59 out2_60 out2_61 out2_62 out2_63 out2_64 out2_65 out2_66 out2_67 out2_68 out2_69 out2_70 out2_71 out2_72 out2_73 out2_74 out2_75 out2_76 out2_77 out2_78 out2_79 out2_80 out2_81 out2_82 out2_83 output0 output1 output2 output3 output4 output5 output6 output7 output8 output9 layer3




**********Input Test****************

v0 in0 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v1 in1 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v2 in2 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v3 in3 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v4 in4 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v5 in5 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v6 in6 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v7 in7 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v8 in8 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v9 in9 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v10 in10 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v11 in11 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v12 in12 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v13 in13 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v14 in14 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v15 in15 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v16 in16 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v17 in17 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v18 in18 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v19 in19 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v20 in20 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v21 in21 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v22 in22 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v23 in23 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v24 in24 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v25 in25 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v26 in26 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v27 in27 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v28 in28 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v29 in29 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v30 in30 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v31 in31 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v32 in32 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v33 in33 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v34 in34 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v35 in35 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v36 in36 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v37 in37 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v38 in38 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v39 in39 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v40 in40 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v41 in41 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v42 in42 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v43 in43 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v44 in44 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v45 in45 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v46 in46 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v47 in47 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v48 in48 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v49 in49 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v50 in50 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v51 in51 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v52 in52 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v53 in53 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v54 in54 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v55 in55 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v56 in56 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v57 in57 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v58 in58 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v59 in59 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v60 in60 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v61 in61 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v62 in62 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v63 in63 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v64 in64 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v65 in65 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v66 in66 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v67 in67 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v68 in68 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v69 in69 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v70 in70 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v71 in71 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v72 in72 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v73 in73 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v74 in74 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v75 in75 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v76 in76 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v77 in77 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v78 in78 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v79 in79 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v80 in80 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v81 in81 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v82 in82 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v83 in83 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v84 in84 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v85 in85 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v86 in86 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v87 in87 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v88 in88 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v89 in89 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v90 in90 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v91 in91 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v92 in92 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v93 in93 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v94 in94 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v95 in95 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v96 in96 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v97 in97 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v98 in98 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v99 in99 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v100 in100 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v101 in101 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v102 in102 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v103 in103 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v104 in104 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v105 in105 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v106 in106 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v107 in107 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v108 in108 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v109 in109 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v110 in110 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v111 in111 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v112 in112 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v113 in113 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v114 in114 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v115 in115 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v116 in116 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v117 in117 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v118 in118 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v119 in119 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v120 in120 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v121 in121 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v122 in122 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v123 in123 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v124 in124 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v125 in125 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v126 in126 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v127 in127 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v128 in128 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v129 in129 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v130 in130 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v131 in131 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v132 in132 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v133 in133 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v134 in134 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v135 in135 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v136 in136 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v137 in137 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v138 in138 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v139 in139 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v140 in140 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v141 in141 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v142 in142 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v143 in143 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v144 in144 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v145 in145 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v146 in146 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v147 in147 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v148 in148 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v149 in149 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v150 in150 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v151 in151 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v152 in152 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v153 in153 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v154 in154 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v155 in155 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v156 in156 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v157 in157 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v158 in158 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v159 in159 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v160 in160 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v161 in161 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v162 in162 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v163 in163 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v164 in164 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v165 in165 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v166 in166 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v167 in167 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v168 in168 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v169 in169 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v170 in170 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v171 in171 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v172 in172 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v173 in173 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v174 in174 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v175 in175 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v176 in176 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v177 in177 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v178 in178 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v179 in179 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v180 in180 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v181 in181 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v182 in182 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v183 in183 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v184 in184 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v185 in185 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v186 in186 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v187 in187 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v188 in188 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v189 in189 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v190 in190 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v191 in191 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v192 in192 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v193 in193 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v194 in194 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v195 in195 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v196 in196 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v197 in197 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v198 in198 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v199 in199 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v200 in200 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v201 in201 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v202 in202 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v203 in203 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v204 in204 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v205 in205 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v206 in206 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v207 in207 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v208 in208 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v209 in209 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v210 in210 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v211 in211 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v212 in212 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v213 in213 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v214 in214 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v215 in215 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v216 in216 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v217 in217 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v218 in218 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v219 in219 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v220 in220 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v221 in221 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v222 in222 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v223 in223 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v224 in224 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v225 in225 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v226 in226 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v227 in227 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v228 in228 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v229 in229 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v230 in230 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v231 in231 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v232 in232 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v233 in233 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v234 in234 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v235 in235 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v236 in236 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v237 in237 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v238 in238 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v239 in239 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v240 in240 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v241 in241 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v242 in242 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v243 in243 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v244 in244 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v245 in245 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v246 in246 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v247 in247 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v248 in248 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v249 in249 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v250 in250 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v251 in251 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v252 in252 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v253 in253 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v254 in254 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v255 in255 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v256 in256 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v257 in257 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v258 in258 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v259 in259 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v260 in260 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v261 in261 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v262 in262 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v263 in263 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v264 in264 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v265 in265 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v266 in266 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v267 in267 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v268 in268 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v269 in269 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v270 in270 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v271 in271 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v272 in272 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v273 in273 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v274 in274 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v275 in275 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v276 in276 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v277 in277 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v278 in278 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v279 in279 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v280 in280 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v281 in281 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v282 in282 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v283 in283 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v284 in284 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v285 in285 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v286 in286 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v287 in287 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v288 in288 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v289 in289 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v290 in290 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v291 in291 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v292 in292 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v293 in293 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v294 in294 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v295 in295 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v296 in296 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v297 in297 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v298 in298 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v299 in299 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v300 in300 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v301 in301 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v302 in302 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v303 in303 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v304 in304 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v305 in305 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v306 in306 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v307 in307 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v308 in308 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v309 in309 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v310 in310 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v311 in311 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v312 in312 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v313 in313 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v314 in314 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v315 in315 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v316 in316 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v317 in317 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v318 in318 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v319 in319 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v320 in320 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v321 in321 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v322 in322 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v323 in323 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v324 in324 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v325 in325 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v326 in326 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v327 in327 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v328 in328 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v329 in329 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v330 in330 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v331 in331 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v332 in332 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v333 in333 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v334 in334 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v335 in335 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v336 in336 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v337 in337 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v338 in338 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v339 in339 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v340 in340 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v341 in341 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v342 in342 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v343 in343 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v344 in344 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v345 in345 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v346 in346 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v347 in347 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v348 in348 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v349 in349 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v350 in350 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v351 in351 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v352 in352 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v353 in353 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v354 in354 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v355 in355 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v356 in356 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v357 in357 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v358 in358 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v359 in359 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v360 in360 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v361 in361 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v362 in362 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v363 in363 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v364 in364 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v365 in365 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v366 in366 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v367 in367 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v368 in368 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v369 in369 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v370 in370 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v371 in371 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v372 in372 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v373 in373 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v374 in374 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v375 in375 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v376 in376 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v377 in377 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v378 in378 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v379 in379 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v380 in380 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v381 in381 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v382 in382 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v383 in383 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v384 in384 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v385 in385 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v386 in386 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v387 in387 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v388 in388 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v389 in389 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v390 in390 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v391 in391 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v392 in392 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v393 in393 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v394 in394 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v395 in395 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v396 in396 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )
v397 in397 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v398 in398 0 PWL( 0n 0 0.100000n -0.800000 4.000000n -0.800000 4.100000n -0.800000 8.000000n -0.800000 )
v399 in399 0 PWL( 0n 0 0.100000n 0.800000 4.000000n 0.800000 4.100000n 0.800000 8.000000n 0.800000 )



vss vss 0 DC VssVal



vdd vdd 0 DC VddVal
.TRAN 0.1n 2*tsampling
.MEASURE TRAN total_energy0 INTEG 'abs(V(vdd)*I(vdd)) + abs(V(vss)*I(vss))' FROM=0*tsampling TO=1*tsampling
.MEASURE TRAN total_energy1 INTEG 'abs(V(vdd)*I(vdd)) + abs(V(vss)*I(vss))' FROM=1*tsampling TO=2*tsampling
.MEAS TRAN VOUT0_0 FIND v(output0) AT=1*tsampling
.MEAS TRAN VOUT1_0 FIND v(output1) AT=1*tsampling
.MEAS TRAN VOUT2_0 FIND v(output2) AT=1*tsampling
.MEAS TRAN VOUT3_0 FIND v(output3) AT=1*tsampling
.MEAS TRAN VOUT4_0 FIND v(output4) AT=1*tsampling
.MEAS TRAN VOUT5_0 FIND v(output5) AT=1*tsampling
.MEAS TRAN VOUT6_0 FIND v(output6) AT=1*tsampling
.MEAS TRAN VOUT7_0 FIND v(output7) AT=1*tsampling
.MEAS TRAN VOUT8_0 FIND v(output8) AT=1*tsampling
.MEAS TRAN VOUT9_0 FIND v(output9) AT=1*tsampling
.MEAS TRAN VOUT0_1 FIND v(output0) AT=2*tsampling
.MEAS TRAN VOUT1_1 FIND v(output1) AT=2*tsampling
.MEAS TRAN VOUT2_1 FIND v(output2) AT=2*tsampling
.MEAS TRAN VOUT3_1 FIND v(output3) AT=2*tsampling
.MEAS TRAN VOUT4_1 FIND v(output4) AT=2*tsampling
.MEAS TRAN VOUT5_1 FIND v(output5) AT=2*tsampling
.MEAS TRAN VOUT6_1 FIND v(output6) AT=2*tsampling
.MEAS TRAN VOUT7_1 FIND v(output7) AT=2*tsampling
.MEAS TRAN VOUT8_1 FIND v(output8) AT=2*tsampling
.MEAS TRAN VOUT9_1 FIND v(output9) AT=2*tsampling
.end