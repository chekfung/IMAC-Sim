.SUBCKT layer3 vdd vss 0 in1 in2 in3 in4 in5 in6 in7 in8 in9 in10 in11 in12 in13 in14 in15 in16 in17 in18 in19 in20 in21 in22 in23 in24 in25 in26 in27 in28 in29 in30 in31 in32 in33 in34 in35 in36 in37 in38 in39 in40 in41 in42 in43 in44 in45 in46 in47 in48 in49 in50 in51 in52 in53 in54 in55 in56 in57 in58 in59 in60 in61 in62 in63 in64 in65 in66 in67 in68 in69 in70 in71 in72 in73 in74 in75 in76 in77 in78 in79 in80 in81 in82 in83 in84 out1 out2 out3 out4 out5 out6 out7 out8 out9 out10 

**********Positive Weighted Array**********
Rwpos1_1 in1_1 sp1_1 78000.000000
Rwpos1_2 in1_2 sp1_2 202000.000000
Rwpos1_3 in1_3 sp1_3 202000.000000
Rwpos1_4 in1_4 sp1_4 202000.000000
Rwpos1_5 in1_5 sp1_5 78000.000000
Rwpos1_6 in1_6 sp1_6 202000.000000
Rwpos1_7 in1_7 sp1_7 202000.000000
Rwpos1_8 in1_8 sp1_8 202000.000000
Rwpos1_9 in1_9 sp1_9 78000.000000
Rwpos1_10 in1_10 sp1_10 78000.000000
Rwpos2_1 in2_1 sp2_1 202000.000000
Rwpos2_2 in2_2 sp2_2 78000.000000
Rwpos2_3 in2_3 sp2_3 78000.000000
Rwpos2_4 in2_4 sp2_4 202000.000000
Rwpos2_5 in2_5 sp2_5 202000.000000
Rwpos2_6 in2_6 sp2_6 78000.000000
Rwpos2_7 in2_7 sp2_7 78000.000000
Rwpos2_8 in2_8 sp2_8 78000.000000
Rwpos2_9 in2_9 sp2_9 202000.000000
Rwpos2_10 in2_10 sp2_10 202000.000000
Rwpos3_1 in3_1 sp3_1 78000.000000
Rwpos3_2 in3_2 sp3_2 78000.000000
Rwpos3_3 in3_3 sp3_3 78000.000000
Rwpos3_4 in3_4 sp3_4 78000.000000
Rwpos3_5 in3_5 sp3_5 202000.000000
Rwpos3_6 in3_6 sp3_6 202000.000000
Rwpos3_7 in3_7 sp3_7 202000.000000
Rwpos3_8 in3_8 sp3_8 78000.000000
Rwpos3_9 in3_9 sp3_9 78000.000000
Rwpos3_10 in3_10 sp3_10 78000.000000
Rwpos4_1 in4_1 sp4_1 78000.000000
Rwpos4_2 in4_2 sp4_2 202000.000000
Rwpos4_3 in4_3 sp4_3 78000.000000
Rwpos4_4 in4_4 sp4_4 202000.000000
Rwpos4_5 in4_5 sp4_5 78000.000000
Rwpos4_6 in4_6 sp4_6 202000.000000
Rwpos4_7 in4_7 sp4_7 78000.000000
Rwpos4_8 in4_8 sp4_8 78000.000000
Rwpos4_9 in4_9 sp4_9 78000.000000
Rwpos4_10 in4_10 sp4_10 202000.000000
Rwpos5_1 in5_1 sp5_1 78000.000000
Rwpos5_2 in5_2 sp5_2 202000.000000
Rwpos5_3 in5_3 sp5_3 78000.000000
Rwpos5_4 in5_4 sp5_4 78000.000000
Rwpos5_5 in5_5 sp5_5 202000.000000
Rwpos5_6 in5_6 sp5_6 202000.000000
Rwpos5_7 in5_7 sp5_7 78000.000000
Rwpos5_8 in5_8 sp5_8 78000.000000
Rwpos5_9 in5_9 sp5_9 78000.000000
Rwpos5_10 in5_10 sp5_10 202000.000000
Rwpos6_1 in6_1 sp6_1 202000.000000
Rwpos6_2 in6_2 sp6_2 78000.000000
Rwpos6_3 in6_3 sp6_3 78000.000000
Rwpos6_4 in6_4 sp6_4 78000.000000
Rwpos6_5 in6_5 sp6_5 78000.000000
Rwpos6_6 in6_6 sp6_6 78000.000000
Rwpos6_7 in6_7 sp6_7 78000.000000
Rwpos6_8 in6_8 sp6_8 202000.000000
Rwpos6_9 in6_9 sp6_9 202000.000000
Rwpos6_10 in6_10 sp6_10 78000.000000
Rwpos7_1 in7_1 sp7_1 78000.000000
Rwpos7_2 in7_2 sp7_2 78000.000000
Rwpos7_3 in7_3 sp7_3 202000.000000
Rwpos7_4 in7_4 sp7_4 202000.000000
Rwpos7_5 in7_5 sp7_5 78000.000000
Rwpos7_6 in7_6 sp7_6 202000.000000
Rwpos7_7 in7_7 sp7_7 78000.000000
Rwpos7_8 in7_8 sp7_8 78000.000000
Rwpos7_9 in7_9 sp7_9 202000.000000
Rwpos7_10 in7_10 sp7_10 202000.000000
Rwpos8_1 in8_1 sp8_1 202000.000000
Rwpos8_2 in8_2 sp8_2 202000.000000
Rwpos8_3 in8_3 sp8_3 78000.000000
Rwpos8_4 in8_4 sp8_4 202000.000000
Rwpos8_5 in8_5 sp8_5 202000.000000
Rwpos8_6 in8_6 sp8_6 78000.000000
Rwpos8_7 in8_7 sp8_7 78000.000000
Rwpos8_8 in8_8 sp8_8 78000.000000
Rwpos8_9 in8_9 sp8_9 78000.000000
Rwpos8_10 in8_10 sp8_10 78000.000000
Rwpos9_1 in9_1 sp9_1 202000.000000
Rwpos9_2 in9_2 sp9_2 202000.000000
Rwpos9_3 in9_3 sp9_3 78000.000000
Rwpos9_4 in9_4 sp9_4 202000.000000
Rwpos9_5 in9_5 sp9_5 78000.000000
Rwpos9_6 in9_6 sp9_6 78000.000000
Rwpos9_7 in9_7 sp9_7 202000.000000
Rwpos9_8 in9_8 sp9_8 78000.000000
Rwpos9_9 in9_9 sp9_9 78000.000000
Rwpos9_10 in9_10 sp9_10 78000.000000
Rwpos10_1 in10_1 sp10_1 202000.000000
Rwpos10_2 in10_2 sp10_2 78000.000000
Rwpos10_3 in10_3 sp10_3 78000.000000
Rwpos10_4 in10_4 sp10_4 78000.000000
Rwpos10_5 in10_5 sp10_5 78000.000000
Rwpos10_6 in10_6 sp10_6 78000.000000
Rwpos10_7 in10_7 sp10_7 202000.000000
Rwpos10_8 in10_8 sp10_8 202000.000000
Rwpos10_9 in10_9 sp10_9 78000.000000
Rwpos10_10 in10_10 sp10_10 78000.000000
Rwpos11_1 in11_1 sp11_1 78000.000000
Rwpos11_2 in11_2 sp11_2 78000.000000
Rwpos11_3 in11_3 sp11_3 202000.000000
Rwpos11_4 in11_4 sp11_4 78000.000000
Rwpos11_5 in11_5 sp11_5 78000.000000
Rwpos11_6 in11_6 sp11_6 78000.000000
Rwpos11_7 in11_7 sp11_7 202000.000000
Rwpos11_8 in11_8 sp11_8 78000.000000
Rwpos11_9 in11_9 sp11_9 78000.000000
Rwpos11_10 in11_10 sp11_10 202000.000000
Rwpos12_1 in12_1 sp12_1 202000.000000
Rwpos12_2 in12_2 sp12_2 202000.000000
Rwpos12_3 in12_3 sp12_3 78000.000000
Rwpos12_4 in12_4 sp12_4 202000.000000
Rwpos12_5 in12_5 sp12_5 78000.000000
Rwpos12_6 in12_6 sp12_6 78000.000000
Rwpos12_7 in12_7 sp12_7 78000.000000
Rwpos12_8 in12_8 sp12_8 202000.000000
Rwpos12_9 in12_9 sp12_9 78000.000000
Rwpos12_10 in12_10 sp12_10 78000.000000
Rwpos13_1 in13_1 sp13_1 78000.000000
Rwpos13_2 in13_2 sp13_2 202000.000000
Rwpos13_3 in13_3 sp13_3 78000.000000
Rwpos13_4 in13_4 sp13_4 78000.000000
Rwpos13_5 in13_5 sp13_5 202000.000000
Rwpos13_6 in13_6 sp13_6 78000.000000
Rwpos13_7 in13_7 sp13_7 78000.000000
Rwpos13_8 in13_8 sp13_8 202000.000000
Rwpos13_9 in13_9 sp13_9 78000.000000
Rwpos13_10 in13_10 sp13_10 202000.000000
Rwpos14_1 in14_1 sp14_1 202000.000000
Rwpos14_2 in14_2 sp14_2 78000.000000
Rwpos14_3 in14_3 sp14_3 78000.000000
Rwpos14_4 in14_4 sp14_4 78000.000000
Rwpos14_5 in14_5 sp14_5 202000.000000
Rwpos14_6 in14_6 sp14_6 202000.000000
Rwpos14_7 in14_7 sp14_7 78000.000000
Rwpos14_8 in14_8 sp14_8 78000.000000
Rwpos14_9 in14_9 sp14_9 78000.000000
Rwpos14_10 in14_10 sp14_10 78000.000000
Rwpos15_1 in15_1 sp15_1 202000.000000
Rwpos15_2 in15_2 sp15_2 78000.000000
Rwpos15_3 in15_3 sp15_3 202000.000000
Rwpos15_4 in15_4 sp15_4 78000.000000
Rwpos15_5 in15_5 sp15_5 78000.000000
Rwpos15_6 in15_6 sp15_6 202000.000000
Rwpos15_7 in15_7 sp15_7 78000.000000
Rwpos15_8 in15_8 sp15_8 202000.000000
Rwpos15_9 in15_9 sp15_9 78000.000000
Rwpos15_10 in15_10 sp15_10 202000.000000
Rwpos16_1 in16_1 sp16_1 202000.000000
Rwpos16_2 in16_2 sp16_2 202000.000000
Rwpos16_3 in16_3 sp16_3 78000.000000
Rwpos16_4 in16_4 sp16_4 202000.000000
Rwpos16_5 in16_5 sp16_5 78000.000000
Rwpos16_6 in16_6 sp16_6 78000.000000
Rwpos16_7 in16_7 sp16_7 78000.000000
Rwpos16_8 in16_8 sp16_8 78000.000000
Rwpos16_9 in16_9 sp16_9 78000.000000
Rwpos16_10 in16_10 sp16_10 202000.000000
Rwpos17_1 in17_1 sp17_1 202000.000000
Rwpos17_2 in17_2 sp17_2 78000.000000
Rwpos17_3 in17_3 sp17_3 202000.000000
Rwpos17_4 in17_4 sp17_4 78000.000000
Rwpos17_5 in17_5 sp17_5 78000.000000
Rwpos17_6 in17_6 sp17_6 78000.000000
Rwpos17_7 in17_7 sp17_7 202000.000000
Rwpos17_8 in17_8 sp17_8 78000.000000
Rwpos17_9 in17_9 sp17_9 202000.000000
Rwpos17_10 in17_10 sp17_10 78000.000000
Rwpos18_1 in18_1 sp18_1 78000.000000
Rwpos18_2 in18_2 sp18_2 202000.000000
Rwpos18_3 in18_3 sp18_3 78000.000000
Rwpos18_4 in18_4 sp18_4 78000.000000
Rwpos18_5 in18_5 sp18_5 202000.000000
Rwpos18_6 in18_6 sp18_6 78000.000000
Rwpos18_7 in18_7 sp18_7 78000.000000
Rwpos18_8 in18_8 sp18_8 202000.000000
Rwpos18_9 in18_9 sp18_9 78000.000000
Rwpos18_10 in18_10 sp18_10 78000.000000
Rwpos19_1 in19_1 sp19_1 202000.000000
Rwpos19_2 in19_2 sp19_2 78000.000000
Rwpos19_3 in19_3 sp19_3 78000.000000
Rwpos19_4 in19_4 sp19_4 78000.000000
Rwpos19_5 in19_5 sp19_5 78000.000000
Rwpos19_6 in19_6 sp19_6 78000.000000
Rwpos19_7 in19_7 sp19_7 78000.000000
Rwpos19_8 in19_8 sp19_8 202000.000000
Rwpos19_9 in19_9 sp19_9 78000.000000
Rwpos19_10 in19_10 sp19_10 202000.000000
Rwpos20_1 in20_1 sp20_1 78000.000000
Rwpos20_2 in20_2 sp20_2 78000.000000
Rwpos20_3 in20_3 sp20_3 78000.000000
Rwpos20_4 in20_4 sp20_4 78000.000000
Rwpos20_5 in20_5 sp20_5 202000.000000
Rwpos20_6 in20_6 sp20_6 78000.000000
Rwpos20_7 in20_7 sp20_7 78000.000000
Rwpos20_8 in20_8 sp20_8 202000.000000
Rwpos20_9 in20_9 sp20_9 78000.000000
Rwpos20_10 in20_10 sp20_10 202000.000000
Rwpos21_1 in21_1 sp21_1 202000.000000
Rwpos21_2 in21_2 sp21_2 202000.000000
Rwpos21_3 in21_3 sp21_3 78000.000000
Rwpos21_4 in21_4 sp21_4 78000.000000
Rwpos21_5 in21_5 sp21_5 78000.000000
Rwpos21_6 in21_6 sp21_6 78000.000000
Rwpos21_7 in21_7 sp21_7 78000.000000
Rwpos21_8 in21_8 sp21_8 78000.000000
Rwpos21_9 in21_9 sp21_9 78000.000000
Rwpos21_10 in21_10 sp21_10 78000.000000
Rwpos22_1 in22_1 sp22_1 202000.000000
Rwpos22_2 in22_2 sp22_2 202000.000000
Rwpos22_3 in22_3 sp22_3 78000.000000
Rwpos22_4 in22_4 sp22_4 78000.000000
Rwpos22_5 in22_5 sp22_5 78000.000000
Rwpos22_6 in22_6 sp22_6 78000.000000
Rwpos22_7 in22_7 sp22_7 202000.000000
Rwpos22_8 in22_8 sp22_8 78000.000000
Rwpos22_9 in22_9 sp22_9 78000.000000
Rwpos22_10 in22_10 sp22_10 78000.000000
Rwpos23_1 in23_1 sp23_1 202000.000000
Rwpos23_2 in23_2 sp23_2 78000.000000
Rwpos23_3 in23_3 sp23_3 202000.000000
Rwpos23_4 in23_4 sp23_4 78000.000000
Rwpos23_5 in23_5 sp23_5 202000.000000
Rwpos23_6 in23_6 sp23_6 78000.000000
Rwpos23_7 in23_7 sp23_7 78000.000000
Rwpos23_8 in23_8 sp23_8 78000.000000
Rwpos23_9 in23_9 sp23_9 78000.000000
Rwpos23_10 in23_10 sp23_10 78000.000000
Rwpos24_1 in24_1 sp24_1 78000.000000
Rwpos24_2 in24_2 sp24_2 78000.000000
Rwpos24_3 in24_3 sp24_3 78000.000000
Rwpos24_4 in24_4 sp24_4 78000.000000
Rwpos24_5 in24_5 sp24_5 78000.000000
Rwpos24_6 in24_6 sp24_6 78000.000000
Rwpos24_7 in24_7 sp24_7 202000.000000
Rwpos24_8 in24_8 sp24_8 202000.000000
Rwpos24_9 in24_9 sp24_9 202000.000000
Rwpos24_10 in24_10 sp24_10 78000.000000
Rwpos25_1 in25_1 sp25_1 202000.000000
Rwpos25_2 in25_2 sp25_2 78000.000000
Rwpos25_3 in25_3 sp25_3 78000.000000
Rwpos25_4 in25_4 sp25_4 78000.000000
Rwpos25_5 in25_5 sp25_5 78000.000000
Rwpos25_6 in25_6 sp25_6 202000.000000
Rwpos25_7 in25_7 sp25_7 78000.000000
Rwpos25_8 in25_8 sp25_8 78000.000000
Rwpos25_9 in25_9 sp25_9 202000.000000
Rwpos25_10 in25_10 sp25_10 78000.000000
Rwpos26_1 in26_1 sp26_1 78000.000000
Rwpos26_2 in26_2 sp26_2 78000.000000
Rwpos26_3 in26_3 sp26_3 202000.000000
Rwpos26_4 in26_4 sp26_4 78000.000000
Rwpos26_5 in26_5 sp26_5 202000.000000
Rwpos26_6 in26_6 sp26_6 202000.000000
Rwpos26_7 in26_7 sp26_7 78000.000000
Rwpos26_8 in26_8 sp26_8 78000.000000
Rwpos26_9 in26_9 sp26_9 78000.000000
Rwpos26_10 in26_10 sp26_10 78000.000000
Rwpos27_1 in27_1 sp27_1 202000.000000
Rwpos27_2 in27_2 sp27_2 202000.000000
Rwpos27_3 in27_3 sp27_3 78000.000000
Rwpos27_4 in27_4 sp27_4 78000.000000
Rwpos27_5 in27_5 sp27_5 78000.000000
Rwpos27_6 in27_6 sp27_6 202000.000000
Rwpos27_7 in27_7 sp27_7 78000.000000
Rwpos27_8 in27_8 sp27_8 78000.000000
Rwpos27_9 in27_9 sp27_9 78000.000000
Rwpos27_10 in27_10 sp27_10 78000.000000
Rwpos28_1 in28_1 sp28_1 78000.000000
Rwpos28_2 in28_2 sp28_2 202000.000000
Rwpos28_3 in28_3 sp28_3 78000.000000
Rwpos28_4 in28_4 sp28_4 78000.000000
Rwpos28_5 in28_5 sp28_5 78000.000000
Rwpos28_6 in28_6 sp28_6 78000.000000
Rwpos28_7 in28_7 sp28_7 78000.000000
Rwpos28_8 in28_8 sp28_8 202000.000000
Rwpos28_9 in28_9 sp28_9 78000.000000
Rwpos28_10 in28_10 sp28_10 202000.000000
Rwpos29_1 in29_1 sp29_1 78000.000000
Rwpos29_2 in29_2 sp29_2 78000.000000
Rwpos29_3 in29_3 sp29_3 78000.000000
Rwpos29_4 in29_4 sp29_4 78000.000000
Rwpos29_5 in29_5 sp29_5 202000.000000
Rwpos29_6 in29_6 sp29_6 78000.000000
Rwpos29_7 in29_7 sp29_7 78000.000000
Rwpos29_8 in29_8 sp29_8 78000.000000
Rwpos29_9 in29_9 sp29_9 202000.000000
Rwpos29_10 in29_10 sp29_10 78000.000000
Rwpos30_1 in30_1 sp30_1 78000.000000
Rwpos30_2 in30_2 sp30_2 202000.000000
Rwpos30_3 in30_3 sp30_3 202000.000000
Rwpos30_4 in30_4 sp30_4 202000.000000
Rwpos30_5 in30_5 sp30_5 78000.000000
Rwpos30_6 in30_6 sp30_6 202000.000000
Rwpos30_7 in30_7 sp30_7 78000.000000
Rwpos30_8 in30_8 sp30_8 202000.000000
Rwpos30_9 in30_9 sp30_9 78000.000000
Rwpos30_10 in30_10 sp30_10 78000.000000
Rwpos31_1 in31_1 sp31_1 202000.000000
Rwpos31_2 in31_2 sp31_2 202000.000000
Rwpos31_3 in31_3 sp31_3 202000.000000
Rwpos31_4 in31_4 sp31_4 78000.000000
Rwpos31_5 in31_5 sp31_5 78000.000000
Rwpos31_6 in31_6 sp31_6 202000.000000
Rwpos31_7 in31_7 sp31_7 202000.000000
Rwpos31_8 in31_8 sp31_8 78000.000000
Rwpos31_9 in31_9 sp31_9 78000.000000
Rwpos31_10 in31_10 sp31_10 78000.000000
Rwpos32_1 in32_1 sp32_1 202000.000000
Rwpos32_2 in32_2 sp32_2 78000.000000
Rwpos32_3 in32_3 sp32_3 202000.000000
Rwpos32_4 in32_4 sp32_4 78000.000000
Rwpos32_5 in32_5 sp32_5 78000.000000
Rwpos32_6 in32_6 sp32_6 78000.000000
Rwpos32_7 in32_7 sp32_7 78000.000000
Rwpos32_8 in32_8 sp32_8 202000.000000
Rwpos32_9 in32_9 sp32_9 78000.000000
Rwpos32_10 in32_10 sp32_10 78000.000000
Rwpos33_1 in33_1 sp33_1 78000.000000
Rwpos33_2 in33_2 sp33_2 78000.000000
Rwpos33_3 in33_3 sp33_3 78000.000000
Rwpos33_4 in33_4 sp33_4 78000.000000
Rwpos33_5 in33_5 sp33_5 202000.000000
Rwpos33_6 in33_6 sp33_6 78000.000000
Rwpos33_7 in33_7 sp33_7 202000.000000
Rwpos33_8 in33_8 sp33_8 78000.000000
Rwpos33_9 in33_9 sp33_9 78000.000000
Rwpos33_10 in33_10 sp33_10 202000.000000
Rwpos34_1 in34_1 sp34_1 202000.000000
Rwpos34_2 in34_2 sp34_2 78000.000000
Rwpos34_3 in34_3 sp34_3 202000.000000
Rwpos34_4 in34_4 sp34_4 202000.000000
Rwpos34_5 in34_5 sp34_5 78000.000000
Rwpos34_6 in34_6 sp34_6 202000.000000
Rwpos34_7 in34_7 sp34_7 78000.000000
Rwpos34_8 in34_8 sp34_8 202000.000000
Rwpos34_9 in34_9 sp34_9 78000.000000
Rwpos34_10 in34_10 sp34_10 78000.000000
Rwpos35_1 in35_1 sp35_1 78000.000000
Rwpos35_2 in35_2 sp35_2 202000.000000
Rwpos35_3 in35_3 sp35_3 78000.000000
Rwpos35_4 in35_4 sp35_4 78000.000000
Rwpos35_5 in35_5 sp35_5 202000.000000
Rwpos35_6 in35_6 sp35_6 202000.000000
Rwpos35_7 in35_7 sp35_7 202000.000000
Rwpos35_8 in35_8 sp35_8 202000.000000
Rwpos35_9 in35_9 sp35_9 78000.000000
Rwpos35_10 in35_10 sp35_10 78000.000000
Rwpos36_1 in36_1 sp36_1 78000.000000
Rwpos36_2 in36_2 sp36_2 78000.000000
Rwpos36_3 in36_3 sp36_3 78000.000000
Rwpos36_4 in36_4 sp36_4 202000.000000
Rwpos36_5 in36_5 sp36_5 78000.000000
Rwpos36_6 in36_6 sp36_6 202000.000000
Rwpos36_7 in36_7 sp36_7 78000.000000
Rwpos36_8 in36_8 sp36_8 202000.000000
Rwpos36_9 in36_9 sp36_9 202000.000000
Rwpos36_10 in36_10 sp36_10 78000.000000
Rwpos37_1 in37_1 sp37_1 78000.000000
Rwpos37_2 in37_2 sp37_2 78000.000000
Rwpos37_3 in37_3 sp37_3 202000.000000
Rwpos37_4 in37_4 sp37_4 202000.000000
Rwpos37_5 in37_5 sp37_5 78000.000000
Rwpos37_6 in37_6 sp37_6 78000.000000
Rwpos37_7 in37_7 sp37_7 78000.000000
Rwpos37_8 in37_8 sp37_8 78000.000000
Rwpos37_9 in37_9 sp37_9 78000.000000
Rwpos37_10 in37_10 sp37_10 202000.000000
Rwpos38_1 in38_1 sp38_1 202000.000000
Rwpos38_2 in38_2 sp38_2 78000.000000
Rwpos38_3 in38_3 sp38_3 78000.000000
Rwpos38_4 in38_4 sp38_4 78000.000000
Rwpos38_5 in38_5 sp38_5 78000.000000
Rwpos38_6 in38_6 sp38_6 202000.000000
Rwpos38_7 in38_7 sp38_7 78000.000000
Rwpos38_8 in38_8 sp38_8 202000.000000
Rwpos38_9 in38_9 sp38_9 78000.000000
Rwpos38_10 in38_10 sp38_10 202000.000000
Rwpos39_1 in39_1 sp39_1 78000.000000
Rwpos39_2 in39_2 sp39_2 202000.000000
Rwpos39_3 in39_3 sp39_3 78000.000000
Rwpos39_4 in39_4 sp39_4 78000.000000
Rwpos39_5 in39_5 sp39_5 78000.000000
Rwpos39_6 in39_6 sp39_6 202000.000000
Rwpos39_7 in39_7 sp39_7 78000.000000
Rwpos39_8 in39_8 sp39_8 202000.000000
Rwpos39_9 in39_9 sp39_9 202000.000000
Rwpos39_10 in39_10 sp39_10 78000.000000
Rwpos40_1 in40_1 sp40_1 202000.000000
Rwpos40_2 in40_2 sp40_2 78000.000000
Rwpos40_3 in40_3 sp40_3 202000.000000
Rwpos40_4 in40_4 sp40_4 78000.000000
Rwpos40_5 in40_5 sp40_5 78000.000000
Rwpos40_6 in40_6 sp40_6 78000.000000
Rwpos40_7 in40_7 sp40_7 78000.000000
Rwpos40_8 in40_8 sp40_8 202000.000000
Rwpos40_9 in40_9 sp40_9 78000.000000
Rwpos40_10 in40_10 sp40_10 202000.000000
Rwpos41_1 in41_1 sp41_1 78000.000000
Rwpos41_2 in41_2 sp41_2 78000.000000
Rwpos41_3 in41_3 sp41_3 78000.000000
Rwpos41_4 in41_4 sp41_4 78000.000000
Rwpos41_5 in41_5 sp41_5 202000.000000
Rwpos41_6 in41_6 sp41_6 78000.000000
Rwpos41_7 in41_7 sp41_7 202000.000000
Rwpos41_8 in41_8 sp41_8 78000.000000
Rwpos41_9 in41_9 sp41_9 78000.000000
Rwpos41_10 in41_10 sp41_10 202000.000000
Rwpos42_1 in42_1 sp42_1 78000.000000
Rwpos42_2 in42_2 sp42_2 78000.000000
Rwpos42_3 in42_3 sp42_3 78000.000000
Rwpos42_4 in42_4 sp42_4 202000.000000
Rwpos42_5 in42_5 sp42_5 202000.000000
Rwpos42_6 in42_6 sp42_6 202000.000000
Rwpos42_7 in42_7 sp42_7 78000.000000
Rwpos42_8 in42_8 sp42_8 78000.000000
Rwpos42_9 in42_9 sp42_9 202000.000000
Rwpos42_10 in42_10 sp42_10 202000.000000
Rwpos43_1 in43_1 sp43_1 78000.000000
Rwpos43_2 in43_2 sp43_2 78000.000000
Rwpos43_3 in43_3 sp43_3 78000.000000
Rwpos43_4 in43_4 sp43_4 202000.000000
Rwpos43_5 in43_5 sp43_5 202000.000000
Rwpos43_6 in43_6 sp43_6 78000.000000
Rwpos43_7 in43_7 sp43_7 202000.000000
Rwpos43_8 in43_8 sp43_8 78000.000000
Rwpos43_9 in43_9 sp43_9 78000.000000
Rwpos43_10 in43_10 sp43_10 202000.000000
Rwpos44_1 in44_1 sp44_1 202000.000000
Rwpos44_2 in44_2 sp44_2 78000.000000
Rwpos44_3 in44_3 sp44_3 78000.000000
Rwpos44_4 in44_4 sp44_4 78000.000000
Rwpos44_5 in44_5 sp44_5 78000.000000
Rwpos44_6 in44_6 sp44_6 78000.000000
Rwpos44_7 in44_7 sp44_7 78000.000000
Rwpos44_8 in44_8 sp44_8 78000.000000
Rwpos44_9 in44_9 sp44_9 202000.000000
Rwpos44_10 in44_10 sp44_10 78000.000000
Rwpos45_1 in45_1 sp45_1 202000.000000
Rwpos45_2 in45_2 sp45_2 78000.000000
Rwpos45_3 in45_3 sp45_3 78000.000000
Rwpos45_4 in45_4 sp45_4 78000.000000
Rwpos45_5 in45_5 sp45_5 202000.000000
Rwpos45_6 in45_6 sp45_6 78000.000000
Rwpos45_7 in45_7 sp45_7 78000.000000
Rwpos45_8 in45_8 sp45_8 202000.000000
Rwpos45_9 in45_9 sp45_9 78000.000000
Rwpos45_10 in45_10 sp45_10 202000.000000
Rwpos46_1 in46_1 sp46_1 78000.000000
Rwpos46_2 in46_2 sp46_2 78000.000000
Rwpos46_3 in46_3 sp46_3 202000.000000
Rwpos46_4 in46_4 sp46_4 78000.000000
Rwpos46_5 in46_5 sp46_5 78000.000000
Rwpos46_6 in46_6 sp46_6 202000.000000
Rwpos46_7 in46_7 sp46_7 78000.000000
Rwpos46_8 in46_8 sp46_8 78000.000000
Rwpos46_9 in46_9 sp46_9 78000.000000
Rwpos46_10 in46_10 sp46_10 78000.000000
Rwpos47_1 in47_1 sp47_1 78000.000000
Rwpos47_2 in47_2 sp47_2 78000.000000
Rwpos47_3 in47_3 sp47_3 78000.000000
Rwpos47_4 in47_4 sp47_4 78000.000000
Rwpos47_5 in47_5 sp47_5 78000.000000
Rwpos47_6 in47_6 sp47_6 202000.000000
Rwpos47_7 in47_7 sp47_7 78000.000000
Rwpos47_8 in47_8 sp47_8 202000.000000
Rwpos47_9 in47_9 sp47_9 202000.000000
Rwpos47_10 in47_10 sp47_10 78000.000000
Rwpos48_1 in48_1 sp48_1 78000.000000
Rwpos48_2 in48_2 sp48_2 78000.000000
Rwpos48_3 in48_3 sp48_3 78000.000000
Rwpos48_4 in48_4 sp48_4 78000.000000
Rwpos48_5 in48_5 sp48_5 78000.000000
Rwpos48_6 in48_6 sp48_6 78000.000000
Rwpos48_7 in48_7 sp48_7 78000.000000
Rwpos48_8 in48_8 sp48_8 78000.000000
Rwpos48_9 in48_9 sp48_9 78000.000000
Rwpos48_10 in48_10 sp48_10 202000.000000
Rwpos49_1 in49_1 sp49_1 202000.000000
Rwpos49_2 in49_2 sp49_2 78000.000000
Rwpos49_3 in49_3 sp49_3 78000.000000
Rwpos49_4 in49_4 sp49_4 202000.000000
Rwpos49_5 in49_5 sp49_5 78000.000000
Rwpos49_6 in49_6 sp49_6 202000.000000
Rwpos49_7 in49_7 sp49_7 78000.000000
Rwpos49_8 in49_8 sp49_8 78000.000000
Rwpos49_9 in49_9 sp49_9 78000.000000
Rwpos49_10 in49_10 sp49_10 202000.000000
Rwpos50_1 in50_1 sp50_1 78000.000000
Rwpos50_2 in50_2 sp50_2 78000.000000
Rwpos50_3 in50_3 sp50_3 78000.000000
Rwpos50_4 in50_4 sp50_4 78000.000000
Rwpos50_5 in50_5 sp50_5 78000.000000
Rwpos50_6 in50_6 sp50_6 202000.000000
Rwpos50_7 in50_7 sp50_7 78000.000000
Rwpos50_8 in50_8 sp50_8 78000.000000
Rwpos50_9 in50_9 sp50_9 78000.000000
Rwpos50_10 in50_10 sp50_10 202000.000000
Rwpos51_1 in51_1 sp51_1 78000.000000
Rwpos51_2 in51_2 sp51_2 202000.000000
Rwpos51_3 in51_3 sp51_3 202000.000000
Rwpos51_4 in51_4 sp51_4 78000.000000
Rwpos51_5 in51_5 sp51_5 78000.000000
Rwpos51_6 in51_6 sp51_6 78000.000000
Rwpos51_7 in51_7 sp51_7 202000.000000
Rwpos51_8 in51_8 sp51_8 78000.000000
Rwpos51_9 in51_9 sp51_9 78000.000000
Rwpos51_10 in51_10 sp51_10 202000.000000
Rwpos52_1 in52_1 sp52_1 202000.000000
Rwpos52_2 in52_2 sp52_2 78000.000000
Rwpos52_3 in52_3 sp52_3 78000.000000
Rwpos52_4 in52_4 sp52_4 202000.000000
Rwpos52_5 in52_5 sp52_5 78000.000000
Rwpos52_6 in52_6 sp52_6 202000.000000
Rwpos52_7 in52_7 sp52_7 78000.000000
Rwpos52_8 in52_8 sp52_8 78000.000000
Rwpos52_9 in52_9 sp52_9 78000.000000
Rwpos52_10 in52_10 sp52_10 202000.000000
Rwpos53_1 in53_1 sp53_1 78000.000000
Rwpos53_2 in53_2 sp53_2 78000.000000
Rwpos53_3 in53_3 sp53_3 78000.000000
Rwpos53_4 in53_4 sp53_4 78000.000000
Rwpos53_5 in53_5 sp53_5 78000.000000
Rwpos53_6 in53_6 sp53_6 78000.000000
Rwpos53_7 in53_7 sp53_7 78000.000000
Rwpos53_8 in53_8 sp53_8 78000.000000
Rwpos53_9 in53_9 sp53_9 78000.000000
Rwpos53_10 in53_10 sp53_10 78000.000000
Rwpos54_1 in54_1 sp54_1 78000.000000
Rwpos54_2 in54_2 sp54_2 202000.000000
Rwpos54_3 in54_3 sp54_3 78000.000000
Rwpos54_4 in54_4 sp54_4 78000.000000
Rwpos54_5 in54_5 sp54_5 78000.000000
Rwpos54_6 in54_6 sp54_6 78000.000000
Rwpos54_7 in54_7 sp54_7 78000.000000
Rwpos54_8 in54_8 sp54_8 78000.000000
Rwpos54_9 in54_9 sp54_9 78000.000000
Rwpos54_10 in54_10 sp54_10 202000.000000
Rwpos55_1 in55_1 sp55_1 78000.000000
Rwpos55_2 in55_2 sp55_2 202000.000000
Rwpos55_3 in55_3 sp55_3 202000.000000
Rwpos55_4 in55_4 sp55_4 78000.000000
Rwpos55_5 in55_5 sp55_5 78000.000000
Rwpos55_6 in55_6 sp55_6 78000.000000
Rwpos55_7 in55_7 sp55_7 202000.000000
Rwpos55_8 in55_8 sp55_8 78000.000000
Rwpos55_9 in55_9 sp55_9 202000.000000
Rwpos55_10 in55_10 sp55_10 78000.000000
Rwpos56_1 in56_1 sp56_1 78000.000000
Rwpos56_2 in56_2 sp56_2 78000.000000
Rwpos56_3 in56_3 sp56_3 202000.000000
Rwpos56_4 in56_4 sp56_4 202000.000000
Rwpos56_5 in56_5 sp56_5 202000.000000
Rwpos56_6 in56_6 sp56_6 78000.000000
Rwpos56_7 in56_7 sp56_7 78000.000000
Rwpos56_8 in56_8 sp56_8 202000.000000
Rwpos56_9 in56_9 sp56_9 78000.000000
Rwpos56_10 in56_10 sp56_10 78000.000000
Rwpos57_1 in57_1 sp57_1 78000.000000
Rwpos57_2 in57_2 sp57_2 78000.000000
Rwpos57_3 in57_3 sp57_3 78000.000000
Rwpos57_4 in57_4 sp57_4 202000.000000
Rwpos57_5 in57_5 sp57_5 78000.000000
Rwpos57_6 in57_6 sp57_6 78000.000000
Rwpos57_7 in57_7 sp57_7 202000.000000
Rwpos57_8 in57_8 sp57_8 202000.000000
Rwpos57_9 in57_9 sp57_9 78000.000000
Rwpos57_10 in57_10 sp57_10 78000.000000
Rwpos58_1 in58_1 sp58_1 202000.000000
Rwpos58_2 in58_2 sp58_2 78000.000000
Rwpos58_3 in58_3 sp58_3 202000.000000
Rwpos58_4 in58_4 sp58_4 78000.000000
Rwpos58_5 in58_5 sp58_5 202000.000000
Rwpos58_6 in58_6 sp58_6 78000.000000
Rwpos58_7 in58_7 sp58_7 78000.000000
Rwpos58_8 in58_8 sp58_8 78000.000000
Rwpos58_9 in58_9 sp58_9 78000.000000
Rwpos58_10 in58_10 sp58_10 78000.000000
Rwpos59_1 in59_1 sp59_1 78000.000000
Rwpos59_2 in59_2 sp59_2 78000.000000
Rwpos59_3 in59_3 sp59_3 78000.000000
Rwpos59_4 in59_4 sp59_4 78000.000000
Rwpos59_5 in59_5 sp59_5 202000.000000
Rwpos59_6 in59_6 sp59_6 202000.000000
Rwpos59_7 in59_7 sp59_7 202000.000000
Rwpos59_8 in59_8 sp59_8 202000.000000
Rwpos59_9 in59_9 sp59_9 202000.000000
Rwpos59_10 in59_10 sp59_10 78000.000000
Rwpos60_1 in60_1 sp60_1 78000.000000
Rwpos60_2 in60_2 sp60_2 78000.000000
Rwpos60_3 in60_3 sp60_3 78000.000000
Rwpos60_4 in60_4 sp60_4 202000.000000
Rwpos60_5 in60_5 sp60_5 78000.000000
Rwpos60_6 in60_6 sp60_6 78000.000000
Rwpos60_7 in60_7 sp60_7 78000.000000
Rwpos60_8 in60_8 sp60_8 78000.000000
Rwpos60_9 in60_9 sp60_9 202000.000000
Rwpos60_10 in60_10 sp60_10 78000.000000
Rwpos61_1 in61_1 sp61_1 202000.000000
Rwpos61_2 in61_2 sp61_2 78000.000000
Rwpos61_3 in61_3 sp61_3 78000.000000
Rwpos61_4 in61_4 sp61_4 202000.000000
Rwpos61_5 in61_5 sp61_5 202000.000000
Rwpos61_6 in61_6 sp61_6 78000.000000
Rwpos61_7 in61_7 sp61_7 202000.000000
Rwpos61_8 in61_8 sp61_8 78000.000000
Rwpos61_9 in61_9 sp61_9 78000.000000
Rwpos61_10 in61_10 sp61_10 78000.000000
Rwpos62_1 in62_1 sp62_1 78000.000000
Rwpos62_2 in62_2 sp62_2 202000.000000
Rwpos62_3 in62_3 sp62_3 202000.000000
Rwpos62_4 in62_4 sp62_4 78000.000000
Rwpos62_5 in62_5 sp62_5 78000.000000
Rwpos62_6 in62_6 sp62_6 78000.000000
Rwpos62_7 in62_7 sp62_7 78000.000000
Rwpos62_8 in62_8 sp62_8 78000.000000
Rwpos62_9 in62_9 sp62_9 202000.000000
Rwpos62_10 in62_10 sp62_10 78000.000000
Rwpos63_1 in63_1 sp63_1 78000.000000
Rwpos63_2 in63_2 sp63_2 78000.000000
Rwpos63_3 in63_3 sp63_3 78000.000000
Rwpos63_4 in63_4 sp63_4 202000.000000
Rwpos63_5 in63_5 sp63_5 202000.000000
Rwpos63_6 in63_6 sp63_6 78000.000000
Rwpos63_7 in63_7 sp63_7 78000.000000
Rwpos63_8 in63_8 sp63_8 202000.000000
Rwpos63_9 in63_9 sp63_9 78000.000000
Rwpos63_10 in63_10 sp63_10 78000.000000
Rwpos64_1 in64_1 sp64_1 78000.000000
Rwpos64_2 in64_2 sp64_2 78000.000000
Rwpos64_3 in64_3 sp64_3 78000.000000
Rwpos64_4 in64_4 sp64_4 78000.000000
Rwpos64_5 in64_5 sp64_5 78000.000000
Rwpos64_6 in64_6 sp64_6 78000.000000
Rwpos64_7 in64_7 sp64_7 78000.000000
Rwpos64_8 in64_8 sp64_8 78000.000000
Rwpos64_9 in64_9 sp64_9 78000.000000
Rwpos64_10 in64_10 sp64_10 78000.000000
Rwpos65_1 in65_1 sp65_1 78000.000000
Rwpos65_2 in65_2 sp65_2 78000.000000
Rwpos65_3 in65_3 sp65_3 202000.000000
Rwpos65_4 in65_4 sp65_4 78000.000000
Rwpos65_5 in65_5 sp65_5 78000.000000
Rwpos65_6 in65_6 sp65_6 78000.000000
Rwpos65_7 in65_7 sp65_7 78000.000000
Rwpos65_8 in65_8 sp65_8 202000.000000
Rwpos65_9 in65_9 sp65_9 202000.000000
Rwpos65_10 in65_10 sp65_10 78000.000000
Rwpos66_1 in66_1 sp66_1 202000.000000
Rwpos66_2 in66_2 sp66_2 202000.000000
Rwpos66_3 in66_3 sp66_3 78000.000000
Rwpos66_4 in66_4 sp66_4 202000.000000
Rwpos66_5 in66_5 sp66_5 78000.000000
Rwpos66_6 in66_6 sp66_6 78000.000000
Rwpos66_7 in66_7 sp66_7 78000.000000
Rwpos66_8 in66_8 sp66_8 78000.000000
Rwpos66_9 in66_9 sp66_9 78000.000000
Rwpos66_10 in66_10 sp66_10 202000.000000
Rwpos67_1 in67_1 sp67_1 202000.000000
Rwpos67_2 in67_2 sp67_2 78000.000000
Rwpos67_3 in67_3 sp67_3 78000.000000
Rwpos67_4 in67_4 sp67_4 78000.000000
Rwpos67_5 in67_5 sp67_5 78000.000000
Rwpos67_6 in67_6 sp67_6 202000.000000
Rwpos67_7 in67_7 sp67_7 78000.000000
Rwpos67_8 in67_8 sp67_8 202000.000000
Rwpos67_9 in67_9 sp67_9 78000.000000
Rwpos67_10 in67_10 sp67_10 78000.000000
Rwpos68_1 in68_1 sp68_1 202000.000000
Rwpos68_2 in68_2 sp68_2 202000.000000
Rwpos68_3 in68_3 sp68_3 78000.000000
Rwpos68_4 in68_4 sp68_4 202000.000000
Rwpos68_5 in68_5 sp68_5 78000.000000
Rwpos68_6 in68_6 sp68_6 78000.000000
Rwpos68_7 in68_7 sp68_7 78000.000000
Rwpos68_8 in68_8 sp68_8 202000.000000
Rwpos68_9 in68_9 sp68_9 202000.000000
Rwpos68_10 in68_10 sp68_10 78000.000000
Rwpos69_1 in69_1 sp69_1 78000.000000
Rwpos69_2 in69_2 sp69_2 202000.000000
Rwpos69_3 in69_3 sp69_3 202000.000000
Rwpos69_4 in69_4 sp69_4 202000.000000
Rwpos69_5 in69_5 sp69_5 78000.000000
Rwpos69_6 in69_6 sp69_6 78000.000000
Rwpos69_7 in69_7 sp69_7 202000.000000
Rwpos69_8 in69_8 sp69_8 202000.000000
Rwpos69_9 in69_9 sp69_9 78000.000000
Rwpos69_10 in69_10 sp69_10 78000.000000
Rwpos70_1 in70_1 sp70_1 78000.000000
Rwpos70_2 in70_2 sp70_2 202000.000000
Rwpos70_3 in70_3 sp70_3 202000.000000
Rwpos70_4 in70_4 sp70_4 78000.000000
Rwpos70_5 in70_5 sp70_5 78000.000000
Rwpos70_6 in70_6 sp70_6 78000.000000
Rwpos70_7 in70_7 sp70_7 202000.000000
Rwpos70_8 in70_8 sp70_8 78000.000000
Rwpos70_9 in70_9 sp70_9 78000.000000
Rwpos70_10 in70_10 sp70_10 202000.000000
Rwpos71_1 in71_1 sp71_1 78000.000000
Rwpos71_2 in71_2 sp71_2 78000.000000
Rwpos71_3 in71_3 sp71_3 202000.000000
Rwpos71_4 in71_4 sp71_4 202000.000000
Rwpos71_5 in71_5 sp71_5 202000.000000
Rwpos71_6 in71_6 sp71_6 78000.000000
Rwpos71_7 in71_7 sp71_7 78000.000000
Rwpos71_8 in71_8 sp71_8 202000.000000
Rwpos71_9 in71_9 sp71_9 78000.000000
Rwpos71_10 in71_10 sp71_10 78000.000000
Rwpos72_1 in72_1 sp72_1 78000.000000
Rwpos72_2 in72_2 sp72_2 78000.000000
Rwpos72_3 in72_3 sp72_3 78000.000000
Rwpos72_4 in72_4 sp72_4 78000.000000
Rwpos72_5 in72_5 sp72_5 78000.000000
Rwpos72_6 in72_6 sp72_6 78000.000000
Rwpos72_7 in72_7 sp72_7 202000.000000
Rwpos72_8 in72_8 sp72_8 78000.000000
Rwpos72_9 in72_9 sp72_9 78000.000000
Rwpos72_10 in72_10 sp72_10 78000.000000
Rwpos73_1 in73_1 sp73_1 202000.000000
Rwpos73_2 in73_2 sp73_2 78000.000000
Rwpos73_3 in73_3 sp73_3 202000.000000
Rwpos73_4 in73_4 sp73_4 202000.000000
Rwpos73_5 in73_5 sp73_5 78000.000000
Rwpos73_6 in73_6 sp73_6 78000.000000
Rwpos73_7 in73_7 sp73_7 202000.000000
Rwpos73_8 in73_8 sp73_8 78000.000000
Rwpos73_9 in73_9 sp73_9 78000.000000
Rwpos73_10 in73_10 sp73_10 78000.000000
Rwpos74_1 in74_1 sp74_1 202000.000000
Rwpos74_2 in74_2 sp74_2 78000.000000
Rwpos74_3 in74_3 sp74_3 78000.000000
Rwpos74_4 in74_4 sp74_4 202000.000000
Rwpos74_5 in74_5 sp74_5 78000.000000
Rwpos74_6 in74_6 sp74_6 202000.000000
Rwpos74_7 in74_7 sp74_7 202000.000000
Rwpos74_8 in74_8 sp74_8 78000.000000
Rwpos74_9 in74_9 sp74_9 78000.000000
Rwpos74_10 in74_10 sp74_10 78000.000000
Rwpos75_1 in75_1 sp75_1 78000.000000
Rwpos75_2 in75_2 sp75_2 78000.000000
Rwpos75_3 in75_3 sp75_3 78000.000000
Rwpos75_4 in75_4 sp75_4 78000.000000
Rwpos75_5 in75_5 sp75_5 202000.000000
Rwpos75_6 in75_6 sp75_6 202000.000000
Rwpos75_7 in75_7 sp75_7 202000.000000
Rwpos75_8 in75_8 sp75_8 202000.000000
Rwpos75_9 in75_9 sp75_9 78000.000000
Rwpos75_10 in75_10 sp75_10 78000.000000
Rwpos76_1 in76_1 sp76_1 78000.000000
Rwpos76_2 in76_2 sp76_2 78000.000000
Rwpos76_3 in76_3 sp76_3 78000.000000
Rwpos76_4 in76_4 sp76_4 202000.000000
Rwpos76_5 in76_5 sp76_5 78000.000000
Rwpos76_6 in76_6 sp76_6 202000.000000
Rwpos76_7 in76_7 sp76_7 78000.000000
Rwpos76_8 in76_8 sp76_8 78000.000000
Rwpos76_9 in76_9 sp76_9 78000.000000
Rwpos76_10 in76_10 sp76_10 78000.000000
Rwpos77_1 in77_1 sp77_1 202000.000000
Rwpos77_2 in77_2 sp77_2 78000.000000
Rwpos77_3 in77_3 sp77_3 202000.000000
Rwpos77_4 in77_4 sp77_4 78000.000000
Rwpos77_5 in77_5 sp77_5 202000.000000
Rwpos77_6 in77_6 sp77_6 78000.000000
Rwpos77_7 in77_7 sp77_7 78000.000000
Rwpos77_8 in77_8 sp77_8 202000.000000
Rwpos77_9 in77_9 sp77_9 78000.000000
Rwpos77_10 in77_10 sp77_10 78000.000000
Rwpos78_1 in78_1 sp78_1 202000.000000
Rwpos78_2 in78_2 sp78_2 202000.000000
Rwpos78_3 in78_3 sp78_3 78000.000000
Rwpos78_4 in78_4 sp78_4 202000.000000
Rwpos78_5 in78_5 sp78_5 202000.000000
Rwpos78_6 in78_6 sp78_6 202000.000000
Rwpos78_7 in78_7 sp78_7 202000.000000
Rwpos78_8 in78_8 sp78_8 78000.000000
Rwpos78_9 in78_9 sp78_9 202000.000000
Rwpos78_10 in78_10 sp78_10 202000.000000
Rwpos79_1 in79_1 sp79_1 78000.000000
Rwpos79_2 in79_2 sp79_2 78000.000000
Rwpos79_3 in79_3 sp79_3 202000.000000
Rwpos79_4 in79_4 sp79_4 202000.000000
Rwpos79_5 in79_5 sp79_5 78000.000000
Rwpos79_6 in79_6 sp79_6 78000.000000
Rwpos79_7 in79_7 sp79_7 78000.000000
Rwpos79_8 in79_8 sp79_8 202000.000000
Rwpos79_9 in79_9 sp79_9 78000.000000
Rwpos79_10 in79_10 sp79_10 78000.000000
Rwpos80_1 in80_1 sp80_1 78000.000000
Rwpos80_2 in80_2 sp80_2 202000.000000
Rwpos80_3 in80_3 sp80_3 202000.000000
Rwpos80_4 in80_4 sp80_4 78000.000000
Rwpos80_5 in80_5 sp80_5 202000.000000
Rwpos80_6 in80_6 sp80_6 78000.000000
Rwpos80_7 in80_7 sp80_7 78000.000000
Rwpos80_8 in80_8 sp80_8 78000.000000
Rwpos80_9 in80_9 sp80_9 78000.000000
Rwpos80_10 in80_10 sp80_10 78000.000000
Rwpos81_1 in81_1 sp81_1 78000.000000
Rwpos81_2 in81_2 sp81_2 78000.000000
Rwpos81_3 in81_3 sp81_3 202000.000000
Rwpos81_4 in81_4 sp81_4 78000.000000
Rwpos81_5 in81_5 sp81_5 202000.000000
Rwpos81_6 in81_6 sp81_6 78000.000000
Rwpos81_7 in81_7 sp81_7 78000.000000
Rwpos81_8 in81_8 sp81_8 78000.000000
Rwpos81_9 in81_9 sp81_9 202000.000000
Rwpos81_10 in81_10 sp81_10 78000.000000
Rwpos82_1 in82_1 sp82_1 78000.000000
Rwpos82_2 in82_2 sp82_2 202000.000000
Rwpos82_3 in82_3 sp82_3 78000.000000
Rwpos82_4 in82_4 sp82_4 202000.000000
Rwpos82_5 in82_5 sp82_5 78000.000000
Rwpos82_6 in82_6 sp82_6 78000.000000
Rwpos82_7 in82_7 sp82_7 78000.000000
Rwpos82_8 in82_8 sp82_8 78000.000000
Rwpos82_9 in82_9 sp82_9 78000.000000
Rwpos82_10 in82_10 sp82_10 78000.000000
Rwpos83_1 in83_1 sp83_1 202000.000000
Rwpos83_2 in83_2 sp83_2 78000.000000
Rwpos83_3 in83_3 sp83_3 78000.000000
Rwpos83_4 in83_4 sp83_4 78000.000000
Rwpos83_5 in83_5 sp83_5 202000.000000
Rwpos83_6 in83_6 sp83_6 202000.000000
Rwpos83_7 in83_7 sp83_7 78000.000000
Rwpos83_8 in83_8 sp83_8 78000.000000
Rwpos83_9 in83_9 sp83_9 78000.000000
Rwpos83_10 in83_10 sp83_10 78000.000000
Rwpos84_1 in84_1 sp84_1 202000.000000
Rwpos84_2 in84_2 sp84_2 78000.000000
Rwpos84_3 in84_3 sp84_3 78000.000000
Rwpos84_4 in84_4 sp84_4 78000.000000
Rwpos84_5 in84_5 sp84_5 202000.000000
Rwpos84_6 in84_6 sp84_6 78000.000000
Rwpos84_7 in84_7 sp84_7 78000.000000
Rwpos84_8 in84_8 sp84_8 78000.000000
Rwpos84_9 in84_9 sp84_9 78000.000000
Rwpos84_10 in84_10 sp84_10 78000.000000


**********Negative Weighted Array**********

Rwneg1_1 in1_1 sn1_1 202000.000000
Rwneg1_2 in1_2 sn1_2 78000.000000
Rwneg1_3 in1_3 sn1_3 78000.000000
Rwneg1_4 in1_4 sn1_4 78000.000000
Rwneg1_5 in1_5 sn1_5 202000.000000
Rwneg1_6 in1_6 sn1_6 78000.000000
Rwneg1_7 in1_7 sn1_7 78000.000000
Rwneg1_8 in1_8 sn1_8 78000.000000
Rwneg1_9 in1_9 sn1_9 202000.000000
Rwneg1_10 in1_10 sn1_10 202000.000000
Rwneg2_1 in2_1 sn2_1 78000.000000
Rwneg2_2 in2_2 sn2_2 202000.000000
Rwneg2_3 in2_3 sn2_3 202000.000000
Rwneg2_4 in2_4 sn2_4 78000.000000
Rwneg2_5 in2_5 sn2_5 78000.000000
Rwneg2_6 in2_6 sn2_6 202000.000000
Rwneg2_7 in2_7 sn2_7 202000.000000
Rwneg2_8 in2_8 sn2_8 202000.000000
Rwneg2_9 in2_9 sn2_9 78000.000000
Rwneg2_10 in2_10 sn2_10 78000.000000
Rwneg3_1 in3_1 sn3_1 202000.000000
Rwneg3_2 in3_2 sn3_2 202000.000000
Rwneg3_3 in3_3 sn3_3 202000.000000
Rwneg3_4 in3_4 sn3_4 202000.000000
Rwneg3_5 in3_5 sn3_5 78000.000000
Rwneg3_6 in3_6 sn3_6 78000.000000
Rwneg3_7 in3_7 sn3_7 78000.000000
Rwneg3_8 in3_8 sn3_8 202000.000000
Rwneg3_9 in3_9 sn3_9 202000.000000
Rwneg3_10 in3_10 sn3_10 202000.000000
Rwneg4_1 in4_1 sn4_1 202000.000000
Rwneg4_2 in4_2 sn4_2 78000.000000
Rwneg4_3 in4_3 sn4_3 202000.000000
Rwneg4_4 in4_4 sn4_4 78000.000000
Rwneg4_5 in4_5 sn4_5 202000.000000
Rwneg4_6 in4_6 sn4_6 78000.000000
Rwneg4_7 in4_7 sn4_7 202000.000000
Rwneg4_8 in4_8 sn4_8 202000.000000
Rwneg4_9 in4_9 sn4_9 202000.000000
Rwneg4_10 in4_10 sn4_10 78000.000000
Rwneg5_1 in5_1 sn5_1 202000.000000
Rwneg5_2 in5_2 sn5_2 78000.000000
Rwneg5_3 in5_3 sn5_3 202000.000000
Rwneg5_4 in5_4 sn5_4 202000.000000
Rwneg5_5 in5_5 sn5_5 78000.000000
Rwneg5_6 in5_6 sn5_6 78000.000000
Rwneg5_7 in5_7 sn5_7 202000.000000
Rwneg5_8 in5_8 sn5_8 202000.000000
Rwneg5_9 in5_9 sn5_9 202000.000000
Rwneg5_10 in5_10 sn5_10 78000.000000
Rwneg6_1 in6_1 sn6_1 78000.000000
Rwneg6_2 in6_2 sn6_2 202000.000000
Rwneg6_3 in6_3 sn6_3 202000.000000
Rwneg6_4 in6_4 sn6_4 202000.000000
Rwneg6_5 in6_5 sn6_5 202000.000000
Rwneg6_6 in6_6 sn6_6 202000.000000
Rwneg6_7 in6_7 sn6_7 202000.000000
Rwneg6_8 in6_8 sn6_8 78000.000000
Rwneg6_9 in6_9 sn6_9 78000.000000
Rwneg6_10 in6_10 sn6_10 202000.000000
Rwneg7_1 in7_1 sn7_1 202000.000000
Rwneg7_2 in7_2 sn7_2 202000.000000
Rwneg7_3 in7_3 sn7_3 78000.000000
Rwneg7_4 in7_4 sn7_4 78000.000000
Rwneg7_5 in7_5 sn7_5 202000.000000
Rwneg7_6 in7_6 sn7_6 78000.000000
Rwneg7_7 in7_7 sn7_7 202000.000000
Rwneg7_8 in7_8 sn7_8 202000.000000
Rwneg7_9 in7_9 sn7_9 78000.000000
Rwneg7_10 in7_10 sn7_10 78000.000000
Rwneg8_1 in8_1 sn8_1 78000.000000
Rwneg8_2 in8_2 sn8_2 78000.000000
Rwneg8_3 in8_3 sn8_3 202000.000000
Rwneg8_4 in8_4 sn8_4 78000.000000
Rwneg8_5 in8_5 sn8_5 78000.000000
Rwneg8_6 in8_6 sn8_6 202000.000000
Rwneg8_7 in8_7 sn8_7 202000.000000
Rwneg8_8 in8_8 sn8_8 202000.000000
Rwneg8_9 in8_9 sn8_9 202000.000000
Rwneg8_10 in8_10 sn8_10 202000.000000
Rwneg9_1 in9_1 sn9_1 78000.000000
Rwneg9_2 in9_2 sn9_2 78000.000000
Rwneg9_3 in9_3 sn9_3 202000.000000
Rwneg9_4 in9_4 sn9_4 78000.000000
Rwneg9_5 in9_5 sn9_5 202000.000000
Rwneg9_6 in9_6 sn9_6 202000.000000
Rwneg9_7 in9_7 sn9_7 78000.000000
Rwneg9_8 in9_8 sn9_8 202000.000000
Rwneg9_9 in9_9 sn9_9 202000.000000
Rwneg9_10 in9_10 sn9_10 202000.000000
Rwneg10_1 in10_1 sn10_1 78000.000000
Rwneg10_2 in10_2 sn10_2 202000.000000
Rwneg10_3 in10_3 sn10_3 202000.000000
Rwneg10_4 in10_4 sn10_4 202000.000000
Rwneg10_5 in10_5 sn10_5 202000.000000
Rwneg10_6 in10_6 sn10_6 202000.000000
Rwneg10_7 in10_7 sn10_7 78000.000000
Rwneg10_8 in10_8 sn10_8 78000.000000
Rwneg10_9 in10_9 sn10_9 202000.000000
Rwneg10_10 in10_10 sn10_10 202000.000000
Rwneg11_1 in11_1 sn11_1 202000.000000
Rwneg11_2 in11_2 sn11_2 202000.000000
Rwneg11_3 in11_3 sn11_3 78000.000000
Rwneg11_4 in11_4 sn11_4 202000.000000
Rwneg11_5 in11_5 sn11_5 202000.000000
Rwneg11_6 in11_6 sn11_6 202000.000000
Rwneg11_7 in11_7 sn11_7 78000.000000
Rwneg11_8 in11_8 sn11_8 202000.000000
Rwneg11_9 in11_9 sn11_9 202000.000000
Rwneg11_10 in11_10 sn11_10 78000.000000
Rwneg12_1 in12_1 sn12_1 78000.000000
Rwneg12_2 in12_2 sn12_2 78000.000000
Rwneg12_3 in12_3 sn12_3 202000.000000
Rwneg12_4 in12_4 sn12_4 78000.000000
Rwneg12_5 in12_5 sn12_5 202000.000000
Rwneg12_6 in12_6 sn12_6 202000.000000
Rwneg12_7 in12_7 sn12_7 202000.000000
Rwneg12_8 in12_8 sn12_8 78000.000000
Rwneg12_9 in12_9 sn12_9 202000.000000
Rwneg12_10 in12_10 sn12_10 202000.000000
Rwneg13_1 in13_1 sn13_1 202000.000000
Rwneg13_2 in13_2 sn13_2 78000.000000
Rwneg13_3 in13_3 sn13_3 202000.000000
Rwneg13_4 in13_4 sn13_4 202000.000000
Rwneg13_5 in13_5 sn13_5 78000.000000
Rwneg13_6 in13_6 sn13_6 202000.000000
Rwneg13_7 in13_7 sn13_7 202000.000000
Rwneg13_8 in13_8 sn13_8 78000.000000
Rwneg13_9 in13_9 sn13_9 202000.000000
Rwneg13_10 in13_10 sn13_10 78000.000000
Rwneg14_1 in14_1 sn14_1 78000.000000
Rwneg14_2 in14_2 sn14_2 202000.000000
Rwneg14_3 in14_3 sn14_3 202000.000000
Rwneg14_4 in14_4 sn14_4 202000.000000
Rwneg14_5 in14_5 sn14_5 78000.000000
Rwneg14_6 in14_6 sn14_6 78000.000000
Rwneg14_7 in14_7 sn14_7 202000.000000
Rwneg14_8 in14_8 sn14_8 202000.000000
Rwneg14_9 in14_9 sn14_9 202000.000000
Rwneg14_10 in14_10 sn14_10 202000.000000
Rwneg15_1 in15_1 sn15_1 78000.000000
Rwneg15_2 in15_2 sn15_2 202000.000000
Rwneg15_3 in15_3 sn15_3 78000.000000
Rwneg15_4 in15_4 sn15_4 202000.000000
Rwneg15_5 in15_5 sn15_5 202000.000000
Rwneg15_6 in15_6 sn15_6 78000.000000
Rwneg15_7 in15_7 sn15_7 202000.000000
Rwneg15_8 in15_8 sn15_8 78000.000000
Rwneg15_9 in15_9 sn15_9 202000.000000
Rwneg15_10 in15_10 sn15_10 78000.000000
Rwneg16_1 in16_1 sn16_1 78000.000000
Rwneg16_2 in16_2 sn16_2 78000.000000
Rwneg16_3 in16_3 sn16_3 202000.000000
Rwneg16_4 in16_4 sn16_4 78000.000000
Rwneg16_5 in16_5 sn16_5 202000.000000
Rwneg16_6 in16_6 sn16_6 202000.000000
Rwneg16_7 in16_7 sn16_7 202000.000000
Rwneg16_8 in16_8 sn16_8 202000.000000
Rwneg16_9 in16_9 sn16_9 202000.000000
Rwneg16_10 in16_10 sn16_10 78000.000000
Rwneg17_1 in17_1 sn17_1 78000.000000
Rwneg17_2 in17_2 sn17_2 202000.000000
Rwneg17_3 in17_3 sn17_3 78000.000000
Rwneg17_4 in17_4 sn17_4 202000.000000
Rwneg17_5 in17_5 sn17_5 202000.000000
Rwneg17_6 in17_6 sn17_6 202000.000000
Rwneg17_7 in17_7 sn17_7 78000.000000
Rwneg17_8 in17_8 sn17_8 202000.000000
Rwneg17_9 in17_9 sn17_9 78000.000000
Rwneg17_10 in17_10 sn17_10 202000.000000
Rwneg18_1 in18_1 sn18_1 202000.000000
Rwneg18_2 in18_2 sn18_2 78000.000000
Rwneg18_3 in18_3 sn18_3 202000.000000
Rwneg18_4 in18_4 sn18_4 202000.000000
Rwneg18_5 in18_5 sn18_5 78000.000000
Rwneg18_6 in18_6 sn18_6 202000.000000
Rwneg18_7 in18_7 sn18_7 202000.000000
Rwneg18_8 in18_8 sn18_8 78000.000000
Rwneg18_9 in18_9 sn18_9 202000.000000
Rwneg18_10 in18_10 sn18_10 202000.000000
Rwneg19_1 in19_1 sn19_1 78000.000000
Rwneg19_2 in19_2 sn19_2 202000.000000
Rwneg19_3 in19_3 sn19_3 202000.000000
Rwneg19_4 in19_4 sn19_4 202000.000000
Rwneg19_5 in19_5 sn19_5 202000.000000
Rwneg19_6 in19_6 sn19_6 202000.000000
Rwneg19_7 in19_7 sn19_7 202000.000000
Rwneg19_8 in19_8 sn19_8 78000.000000
Rwneg19_9 in19_9 sn19_9 202000.000000
Rwneg19_10 in19_10 sn19_10 78000.000000
Rwneg20_1 in20_1 sn20_1 202000.000000
Rwneg20_2 in20_2 sn20_2 202000.000000
Rwneg20_3 in20_3 sn20_3 202000.000000
Rwneg20_4 in20_4 sn20_4 202000.000000
Rwneg20_5 in20_5 sn20_5 78000.000000
Rwneg20_6 in20_6 sn20_6 202000.000000
Rwneg20_7 in20_7 sn20_7 202000.000000
Rwneg20_8 in20_8 sn20_8 78000.000000
Rwneg20_9 in20_9 sn20_9 202000.000000
Rwneg20_10 in20_10 sn20_10 78000.000000
Rwneg21_1 in21_1 sn21_1 78000.000000
Rwneg21_2 in21_2 sn21_2 78000.000000
Rwneg21_3 in21_3 sn21_3 202000.000000
Rwneg21_4 in21_4 sn21_4 202000.000000
Rwneg21_5 in21_5 sn21_5 202000.000000
Rwneg21_6 in21_6 sn21_6 202000.000000
Rwneg21_7 in21_7 sn21_7 202000.000000
Rwneg21_8 in21_8 sn21_8 202000.000000
Rwneg21_9 in21_9 sn21_9 202000.000000
Rwneg21_10 in21_10 sn21_10 202000.000000
Rwneg22_1 in22_1 sn22_1 78000.000000
Rwneg22_2 in22_2 sn22_2 78000.000000
Rwneg22_3 in22_3 sn22_3 202000.000000
Rwneg22_4 in22_4 sn22_4 202000.000000
Rwneg22_5 in22_5 sn22_5 202000.000000
Rwneg22_6 in22_6 sn22_6 202000.000000
Rwneg22_7 in22_7 sn22_7 78000.000000
Rwneg22_8 in22_8 sn22_8 202000.000000
Rwneg22_9 in22_9 sn22_9 202000.000000
Rwneg22_10 in22_10 sn22_10 202000.000000
Rwneg23_1 in23_1 sn23_1 78000.000000
Rwneg23_2 in23_2 sn23_2 202000.000000
Rwneg23_3 in23_3 sn23_3 78000.000000
Rwneg23_4 in23_4 sn23_4 202000.000000
Rwneg23_5 in23_5 sn23_5 78000.000000
Rwneg23_6 in23_6 sn23_6 202000.000000
Rwneg23_7 in23_7 sn23_7 202000.000000
Rwneg23_8 in23_8 sn23_8 202000.000000
Rwneg23_9 in23_9 sn23_9 202000.000000
Rwneg23_10 in23_10 sn23_10 202000.000000
Rwneg24_1 in24_1 sn24_1 202000.000000
Rwneg24_2 in24_2 sn24_2 202000.000000
Rwneg24_3 in24_3 sn24_3 202000.000000
Rwneg24_4 in24_4 sn24_4 202000.000000
Rwneg24_5 in24_5 sn24_5 202000.000000
Rwneg24_6 in24_6 sn24_6 202000.000000
Rwneg24_7 in24_7 sn24_7 78000.000000
Rwneg24_8 in24_8 sn24_8 78000.000000
Rwneg24_9 in24_9 sn24_9 78000.000000
Rwneg24_10 in24_10 sn24_10 202000.000000
Rwneg25_1 in25_1 sn25_1 78000.000000
Rwneg25_2 in25_2 sn25_2 202000.000000
Rwneg25_3 in25_3 sn25_3 202000.000000
Rwneg25_4 in25_4 sn25_4 202000.000000
Rwneg25_5 in25_5 sn25_5 202000.000000
Rwneg25_6 in25_6 sn25_6 78000.000000
Rwneg25_7 in25_7 sn25_7 202000.000000
Rwneg25_8 in25_8 sn25_8 202000.000000
Rwneg25_9 in25_9 sn25_9 78000.000000
Rwneg25_10 in25_10 sn25_10 202000.000000
Rwneg26_1 in26_1 sn26_1 202000.000000
Rwneg26_2 in26_2 sn26_2 202000.000000
Rwneg26_3 in26_3 sn26_3 78000.000000
Rwneg26_4 in26_4 sn26_4 202000.000000
Rwneg26_5 in26_5 sn26_5 78000.000000
Rwneg26_6 in26_6 sn26_6 78000.000000
Rwneg26_7 in26_7 sn26_7 202000.000000
Rwneg26_8 in26_8 sn26_8 202000.000000
Rwneg26_9 in26_9 sn26_9 202000.000000
Rwneg26_10 in26_10 sn26_10 202000.000000
Rwneg27_1 in27_1 sn27_1 78000.000000
Rwneg27_2 in27_2 sn27_2 78000.000000
Rwneg27_3 in27_3 sn27_3 202000.000000
Rwneg27_4 in27_4 sn27_4 202000.000000
Rwneg27_5 in27_5 sn27_5 202000.000000
Rwneg27_6 in27_6 sn27_6 78000.000000
Rwneg27_7 in27_7 sn27_7 202000.000000
Rwneg27_8 in27_8 sn27_8 202000.000000
Rwneg27_9 in27_9 sn27_9 202000.000000
Rwneg27_10 in27_10 sn27_10 202000.000000
Rwneg28_1 in28_1 sn28_1 202000.000000
Rwneg28_2 in28_2 sn28_2 78000.000000
Rwneg28_3 in28_3 sn28_3 202000.000000
Rwneg28_4 in28_4 sn28_4 202000.000000
Rwneg28_5 in28_5 sn28_5 202000.000000
Rwneg28_6 in28_6 sn28_6 202000.000000
Rwneg28_7 in28_7 sn28_7 202000.000000
Rwneg28_8 in28_8 sn28_8 78000.000000
Rwneg28_9 in28_9 sn28_9 202000.000000
Rwneg28_10 in28_10 sn28_10 78000.000000
Rwneg29_1 in29_1 sn29_1 202000.000000
Rwneg29_2 in29_2 sn29_2 202000.000000
Rwneg29_3 in29_3 sn29_3 202000.000000
Rwneg29_4 in29_4 sn29_4 202000.000000
Rwneg29_5 in29_5 sn29_5 78000.000000
Rwneg29_6 in29_6 sn29_6 202000.000000
Rwneg29_7 in29_7 sn29_7 202000.000000
Rwneg29_8 in29_8 sn29_8 202000.000000
Rwneg29_9 in29_9 sn29_9 78000.000000
Rwneg29_10 in29_10 sn29_10 202000.000000
Rwneg30_1 in30_1 sn30_1 202000.000000
Rwneg30_2 in30_2 sn30_2 78000.000000
Rwneg30_3 in30_3 sn30_3 78000.000000
Rwneg30_4 in30_4 sn30_4 78000.000000
Rwneg30_5 in30_5 sn30_5 202000.000000
Rwneg30_6 in30_6 sn30_6 78000.000000
Rwneg30_7 in30_7 sn30_7 202000.000000
Rwneg30_8 in30_8 sn30_8 78000.000000
Rwneg30_9 in30_9 sn30_9 202000.000000
Rwneg30_10 in30_10 sn30_10 202000.000000
Rwneg31_1 in31_1 sn31_1 78000.000000
Rwneg31_2 in31_2 sn31_2 78000.000000
Rwneg31_3 in31_3 sn31_3 78000.000000
Rwneg31_4 in31_4 sn31_4 202000.000000
Rwneg31_5 in31_5 sn31_5 202000.000000
Rwneg31_6 in31_6 sn31_6 78000.000000
Rwneg31_7 in31_7 sn31_7 78000.000000
Rwneg31_8 in31_8 sn31_8 202000.000000
Rwneg31_9 in31_9 sn31_9 202000.000000
Rwneg31_10 in31_10 sn31_10 202000.000000
Rwneg32_1 in32_1 sn32_1 78000.000000
Rwneg32_2 in32_2 sn32_2 202000.000000
Rwneg32_3 in32_3 sn32_3 78000.000000
Rwneg32_4 in32_4 sn32_4 202000.000000
Rwneg32_5 in32_5 sn32_5 202000.000000
Rwneg32_6 in32_6 sn32_6 202000.000000
Rwneg32_7 in32_7 sn32_7 202000.000000
Rwneg32_8 in32_8 sn32_8 78000.000000
Rwneg32_9 in32_9 sn32_9 202000.000000
Rwneg32_10 in32_10 sn32_10 202000.000000
Rwneg33_1 in33_1 sn33_1 202000.000000
Rwneg33_2 in33_2 sn33_2 202000.000000
Rwneg33_3 in33_3 sn33_3 202000.000000
Rwneg33_4 in33_4 sn33_4 202000.000000
Rwneg33_5 in33_5 sn33_5 78000.000000
Rwneg33_6 in33_6 sn33_6 202000.000000
Rwneg33_7 in33_7 sn33_7 78000.000000
Rwneg33_8 in33_8 sn33_8 202000.000000
Rwneg33_9 in33_9 sn33_9 202000.000000
Rwneg33_10 in33_10 sn33_10 78000.000000
Rwneg34_1 in34_1 sn34_1 78000.000000
Rwneg34_2 in34_2 sn34_2 202000.000000
Rwneg34_3 in34_3 sn34_3 78000.000000
Rwneg34_4 in34_4 sn34_4 78000.000000
Rwneg34_5 in34_5 sn34_5 202000.000000
Rwneg34_6 in34_6 sn34_6 78000.000000
Rwneg34_7 in34_7 sn34_7 202000.000000
Rwneg34_8 in34_8 sn34_8 78000.000000
Rwneg34_9 in34_9 sn34_9 202000.000000
Rwneg34_10 in34_10 sn34_10 202000.000000
Rwneg35_1 in35_1 sn35_1 202000.000000
Rwneg35_2 in35_2 sn35_2 78000.000000
Rwneg35_3 in35_3 sn35_3 202000.000000
Rwneg35_4 in35_4 sn35_4 202000.000000
Rwneg35_5 in35_5 sn35_5 78000.000000
Rwneg35_6 in35_6 sn35_6 78000.000000
Rwneg35_7 in35_7 sn35_7 78000.000000
Rwneg35_8 in35_8 sn35_8 78000.000000
Rwneg35_9 in35_9 sn35_9 202000.000000
Rwneg35_10 in35_10 sn35_10 202000.000000
Rwneg36_1 in36_1 sn36_1 202000.000000
Rwneg36_2 in36_2 sn36_2 202000.000000
Rwneg36_3 in36_3 sn36_3 202000.000000
Rwneg36_4 in36_4 sn36_4 78000.000000
Rwneg36_5 in36_5 sn36_5 202000.000000
Rwneg36_6 in36_6 sn36_6 78000.000000
Rwneg36_7 in36_7 sn36_7 202000.000000
Rwneg36_8 in36_8 sn36_8 78000.000000
Rwneg36_9 in36_9 sn36_9 78000.000000
Rwneg36_10 in36_10 sn36_10 202000.000000
Rwneg37_1 in37_1 sn37_1 202000.000000
Rwneg37_2 in37_2 sn37_2 202000.000000
Rwneg37_3 in37_3 sn37_3 78000.000000
Rwneg37_4 in37_4 sn37_4 78000.000000
Rwneg37_5 in37_5 sn37_5 202000.000000
Rwneg37_6 in37_6 sn37_6 202000.000000
Rwneg37_7 in37_7 sn37_7 202000.000000
Rwneg37_8 in37_8 sn37_8 202000.000000
Rwneg37_9 in37_9 sn37_9 202000.000000
Rwneg37_10 in37_10 sn37_10 78000.000000
Rwneg38_1 in38_1 sn38_1 78000.000000
Rwneg38_2 in38_2 sn38_2 202000.000000
Rwneg38_3 in38_3 sn38_3 202000.000000
Rwneg38_4 in38_4 sn38_4 202000.000000
Rwneg38_5 in38_5 sn38_5 202000.000000
Rwneg38_6 in38_6 sn38_6 78000.000000
Rwneg38_7 in38_7 sn38_7 202000.000000
Rwneg38_8 in38_8 sn38_8 78000.000000
Rwneg38_9 in38_9 sn38_9 202000.000000
Rwneg38_10 in38_10 sn38_10 78000.000000
Rwneg39_1 in39_1 sn39_1 202000.000000
Rwneg39_2 in39_2 sn39_2 78000.000000
Rwneg39_3 in39_3 sn39_3 202000.000000
Rwneg39_4 in39_4 sn39_4 202000.000000
Rwneg39_5 in39_5 sn39_5 202000.000000
Rwneg39_6 in39_6 sn39_6 78000.000000
Rwneg39_7 in39_7 sn39_7 202000.000000
Rwneg39_8 in39_8 sn39_8 78000.000000
Rwneg39_9 in39_9 sn39_9 78000.000000
Rwneg39_10 in39_10 sn39_10 202000.000000
Rwneg40_1 in40_1 sn40_1 78000.000000
Rwneg40_2 in40_2 sn40_2 202000.000000
Rwneg40_3 in40_3 sn40_3 78000.000000
Rwneg40_4 in40_4 sn40_4 202000.000000
Rwneg40_5 in40_5 sn40_5 202000.000000
Rwneg40_6 in40_6 sn40_6 202000.000000
Rwneg40_7 in40_7 sn40_7 202000.000000
Rwneg40_8 in40_8 sn40_8 78000.000000
Rwneg40_9 in40_9 sn40_9 202000.000000
Rwneg40_10 in40_10 sn40_10 78000.000000
Rwneg41_1 in41_1 sn41_1 202000.000000
Rwneg41_2 in41_2 sn41_2 202000.000000
Rwneg41_3 in41_3 sn41_3 202000.000000
Rwneg41_4 in41_4 sn41_4 202000.000000
Rwneg41_5 in41_5 sn41_5 78000.000000
Rwneg41_6 in41_6 sn41_6 202000.000000
Rwneg41_7 in41_7 sn41_7 78000.000000
Rwneg41_8 in41_8 sn41_8 202000.000000
Rwneg41_9 in41_9 sn41_9 202000.000000
Rwneg41_10 in41_10 sn41_10 78000.000000
Rwneg42_1 in42_1 sn42_1 202000.000000
Rwneg42_2 in42_2 sn42_2 202000.000000
Rwneg42_3 in42_3 sn42_3 202000.000000
Rwneg42_4 in42_4 sn42_4 78000.000000
Rwneg42_5 in42_5 sn42_5 78000.000000
Rwneg42_6 in42_6 sn42_6 78000.000000
Rwneg42_7 in42_7 sn42_7 202000.000000
Rwneg42_8 in42_8 sn42_8 202000.000000
Rwneg42_9 in42_9 sn42_9 78000.000000
Rwneg42_10 in42_10 sn42_10 78000.000000
Rwneg43_1 in43_1 sn43_1 202000.000000
Rwneg43_2 in43_2 sn43_2 202000.000000
Rwneg43_3 in43_3 sn43_3 202000.000000
Rwneg43_4 in43_4 sn43_4 78000.000000
Rwneg43_5 in43_5 sn43_5 78000.000000
Rwneg43_6 in43_6 sn43_6 202000.000000
Rwneg43_7 in43_7 sn43_7 78000.000000
Rwneg43_8 in43_8 sn43_8 202000.000000
Rwneg43_9 in43_9 sn43_9 202000.000000
Rwneg43_10 in43_10 sn43_10 78000.000000
Rwneg44_1 in44_1 sn44_1 78000.000000
Rwneg44_2 in44_2 sn44_2 202000.000000
Rwneg44_3 in44_3 sn44_3 202000.000000
Rwneg44_4 in44_4 sn44_4 202000.000000
Rwneg44_5 in44_5 sn44_5 202000.000000
Rwneg44_6 in44_6 sn44_6 202000.000000
Rwneg44_7 in44_7 sn44_7 202000.000000
Rwneg44_8 in44_8 sn44_8 202000.000000
Rwneg44_9 in44_9 sn44_9 78000.000000
Rwneg44_10 in44_10 sn44_10 202000.000000
Rwneg45_1 in45_1 sn45_1 78000.000000
Rwneg45_2 in45_2 sn45_2 202000.000000
Rwneg45_3 in45_3 sn45_3 202000.000000
Rwneg45_4 in45_4 sn45_4 202000.000000
Rwneg45_5 in45_5 sn45_5 78000.000000
Rwneg45_6 in45_6 sn45_6 202000.000000
Rwneg45_7 in45_7 sn45_7 202000.000000
Rwneg45_8 in45_8 sn45_8 78000.000000
Rwneg45_9 in45_9 sn45_9 202000.000000
Rwneg45_10 in45_10 sn45_10 78000.000000
Rwneg46_1 in46_1 sn46_1 202000.000000
Rwneg46_2 in46_2 sn46_2 202000.000000
Rwneg46_3 in46_3 sn46_3 78000.000000
Rwneg46_4 in46_4 sn46_4 202000.000000
Rwneg46_5 in46_5 sn46_5 202000.000000
Rwneg46_6 in46_6 sn46_6 78000.000000
Rwneg46_7 in46_7 sn46_7 202000.000000
Rwneg46_8 in46_8 sn46_8 202000.000000
Rwneg46_9 in46_9 sn46_9 202000.000000
Rwneg46_10 in46_10 sn46_10 202000.000000
Rwneg47_1 in47_1 sn47_1 202000.000000
Rwneg47_2 in47_2 sn47_2 202000.000000
Rwneg47_3 in47_3 sn47_3 202000.000000
Rwneg47_4 in47_4 sn47_4 202000.000000
Rwneg47_5 in47_5 sn47_5 202000.000000
Rwneg47_6 in47_6 sn47_6 78000.000000
Rwneg47_7 in47_7 sn47_7 202000.000000
Rwneg47_8 in47_8 sn47_8 78000.000000
Rwneg47_9 in47_9 sn47_9 78000.000000
Rwneg47_10 in47_10 sn47_10 202000.000000
Rwneg48_1 in48_1 sn48_1 202000.000000
Rwneg48_2 in48_2 sn48_2 202000.000000
Rwneg48_3 in48_3 sn48_3 202000.000000
Rwneg48_4 in48_4 sn48_4 202000.000000
Rwneg48_5 in48_5 sn48_5 202000.000000
Rwneg48_6 in48_6 sn48_6 202000.000000
Rwneg48_7 in48_7 sn48_7 202000.000000
Rwneg48_8 in48_8 sn48_8 202000.000000
Rwneg48_9 in48_9 sn48_9 202000.000000
Rwneg48_10 in48_10 sn48_10 78000.000000
Rwneg49_1 in49_1 sn49_1 78000.000000
Rwneg49_2 in49_2 sn49_2 202000.000000
Rwneg49_3 in49_3 sn49_3 202000.000000
Rwneg49_4 in49_4 sn49_4 78000.000000
Rwneg49_5 in49_5 sn49_5 202000.000000
Rwneg49_6 in49_6 sn49_6 78000.000000
Rwneg49_7 in49_7 sn49_7 202000.000000
Rwneg49_8 in49_8 sn49_8 202000.000000
Rwneg49_9 in49_9 sn49_9 202000.000000
Rwneg49_10 in49_10 sn49_10 78000.000000
Rwneg50_1 in50_1 sn50_1 202000.000000
Rwneg50_2 in50_2 sn50_2 202000.000000
Rwneg50_3 in50_3 sn50_3 202000.000000
Rwneg50_4 in50_4 sn50_4 202000.000000
Rwneg50_5 in50_5 sn50_5 202000.000000
Rwneg50_6 in50_6 sn50_6 78000.000000
Rwneg50_7 in50_7 sn50_7 202000.000000
Rwneg50_8 in50_8 sn50_8 202000.000000
Rwneg50_9 in50_9 sn50_9 202000.000000
Rwneg50_10 in50_10 sn50_10 78000.000000
Rwneg51_1 in51_1 sn51_1 202000.000000
Rwneg51_2 in51_2 sn51_2 78000.000000
Rwneg51_3 in51_3 sn51_3 78000.000000
Rwneg51_4 in51_4 sn51_4 202000.000000
Rwneg51_5 in51_5 sn51_5 202000.000000
Rwneg51_6 in51_6 sn51_6 202000.000000
Rwneg51_7 in51_7 sn51_7 78000.000000
Rwneg51_8 in51_8 sn51_8 202000.000000
Rwneg51_9 in51_9 sn51_9 202000.000000
Rwneg51_10 in51_10 sn51_10 78000.000000
Rwneg52_1 in52_1 sn52_1 78000.000000
Rwneg52_2 in52_2 sn52_2 202000.000000
Rwneg52_3 in52_3 sn52_3 202000.000000
Rwneg52_4 in52_4 sn52_4 78000.000000
Rwneg52_5 in52_5 sn52_5 202000.000000
Rwneg52_6 in52_6 sn52_6 78000.000000
Rwneg52_7 in52_7 sn52_7 202000.000000
Rwneg52_8 in52_8 sn52_8 202000.000000
Rwneg52_9 in52_9 sn52_9 202000.000000
Rwneg52_10 in52_10 sn52_10 78000.000000
Rwneg53_1 in53_1 sn53_1 202000.000000
Rwneg53_2 in53_2 sn53_2 202000.000000
Rwneg53_3 in53_3 sn53_3 202000.000000
Rwneg53_4 in53_4 sn53_4 202000.000000
Rwneg53_5 in53_5 sn53_5 202000.000000
Rwneg53_6 in53_6 sn53_6 202000.000000
Rwneg53_7 in53_7 sn53_7 202000.000000
Rwneg53_8 in53_8 sn53_8 202000.000000
Rwneg53_9 in53_9 sn53_9 202000.000000
Rwneg53_10 in53_10 sn53_10 202000.000000
Rwneg54_1 in54_1 sn54_1 202000.000000
Rwneg54_2 in54_2 sn54_2 78000.000000
Rwneg54_3 in54_3 sn54_3 202000.000000
Rwneg54_4 in54_4 sn54_4 202000.000000
Rwneg54_5 in54_5 sn54_5 202000.000000
Rwneg54_6 in54_6 sn54_6 202000.000000
Rwneg54_7 in54_7 sn54_7 202000.000000
Rwneg54_8 in54_8 sn54_8 202000.000000
Rwneg54_9 in54_9 sn54_9 202000.000000
Rwneg54_10 in54_10 sn54_10 78000.000000
Rwneg55_1 in55_1 sn55_1 202000.000000
Rwneg55_2 in55_2 sn55_2 78000.000000
Rwneg55_3 in55_3 sn55_3 78000.000000
Rwneg55_4 in55_4 sn55_4 202000.000000
Rwneg55_5 in55_5 sn55_5 202000.000000
Rwneg55_6 in55_6 sn55_6 202000.000000
Rwneg55_7 in55_7 sn55_7 78000.000000
Rwneg55_8 in55_8 sn55_8 202000.000000
Rwneg55_9 in55_9 sn55_9 78000.000000
Rwneg55_10 in55_10 sn55_10 202000.000000
Rwneg56_1 in56_1 sn56_1 202000.000000
Rwneg56_2 in56_2 sn56_2 202000.000000
Rwneg56_3 in56_3 sn56_3 78000.000000
Rwneg56_4 in56_4 sn56_4 78000.000000
Rwneg56_5 in56_5 sn56_5 78000.000000
Rwneg56_6 in56_6 sn56_6 202000.000000
Rwneg56_7 in56_7 sn56_7 202000.000000
Rwneg56_8 in56_8 sn56_8 78000.000000
Rwneg56_9 in56_9 sn56_9 202000.000000
Rwneg56_10 in56_10 sn56_10 202000.000000
Rwneg57_1 in57_1 sn57_1 202000.000000
Rwneg57_2 in57_2 sn57_2 202000.000000
Rwneg57_3 in57_3 sn57_3 202000.000000
Rwneg57_4 in57_4 sn57_4 78000.000000
Rwneg57_5 in57_5 sn57_5 202000.000000
Rwneg57_6 in57_6 sn57_6 202000.000000
Rwneg57_7 in57_7 sn57_7 78000.000000
Rwneg57_8 in57_8 sn57_8 78000.000000
Rwneg57_9 in57_9 sn57_9 202000.000000
Rwneg57_10 in57_10 sn57_10 202000.000000
Rwneg58_1 in58_1 sn58_1 78000.000000
Rwneg58_2 in58_2 sn58_2 202000.000000
Rwneg58_3 in58_3 sn58_3 78000.000000
Rwneg58_4 in58_4 sn58_4 202000.000000
Rwneg58_5 in58_5 sn58_5 78000.000000
Rwneg58_6 in58_6 sn58_6 202000.000000
Rwneg58_7 in58_7 sn58_7 202000.000000
Rwneg58_8 in58_8 sn58_8 202000.000000
Rwneg58_9 in58_9 sn58_9 202000.000000
Rwneg58_10 in58_10 sn58_10 202000.000000
Rwneg59_1 in59_1 sn59_1 202000.000000
Rwneg59_2 in59_2 sn59_2 202000.000000
Rwneg59_3 in59_3 sn59_3 202000.000000
Rwneg59_4 in59_4 sn59_4 202000.000000
Rwneg59_5 in59_5 sn59_5 78000.000000
Rwneg59_6 in59_6 sn59_6 78000.000000
Rwneg59_7 in59_7 sn59_7 78000.000000
Rwneg59_8 in59_8 sn59_8 78000.000000
Rwneg59_9 in59_9 sn59_9 78000.000000
Rwneg59_10 in59_10 sn59_10 202000.000000
Rwneg60_1 in60_1 sn60_1 202000.000000
Rwneg60_2 in60_2 sn60_2 202000.000000
Rwneg60_3 in60_3 sn60_3 202000.000000
Rwneg60_4 in60_4 sn60_4 78000.000000
Rwneg60_5 in60_5 sn60_5 202000.000000
Rwneg60_6 in60_6 sn60_6 202000.000000
Rwneg60_7 in60_7 sn60_7 202000.000000
Rwneg60_8 in60_8 sn60_8 202000.000000
Rwneg60_9 in60_9 sn60_9 78000.000000
Rwneg60_10 in60_10 sn60_10 202000.000000
Rwneg61_1 in61_1 sn61_1 78000.000000
Rwneg61_2 in61_2 sn61_2 202000.000000
Rwneg61_3 in61_3 sn61_3 202000.000000
Rwneg61_4 in61_4 sn61_4 78000.000000
Rwneg61_5 in61_5 sn61_5 78000.000000
Rwneg61_6 in61_6 sn61_6 202000.000000
Rwneg61_7 in61_7 sn61_7 78000.000000
Rwneg61_8 in61_8 sn61_8 202000.000000
Rwneg61_9 in61_9 sn61_9 202000.000000
Rwneg61_10 in61_10 sn61_10 202000.000000
Rwneg62_1 in62_1 sn62_1 202000.000000
Rwneg62_2 in62_2 sn62_2 78000.000000
Rwneg62_3 in62_3 sn62_3 78000.000000
Rwneg62_4 in62_4 sn62_4 202000.000000
Rwneg62_5 in62_5 sn62_5 202000.000000
Rwneg62_6 in62_6 sn62_6 202000.000000
Rwneg62_7 in62_7 sn62_7 202000.000000
Rwneg62_8 in62_8 sn62_8 202000.000000
Rwneg62_9 in62_9 sn62_9 78000.000000
Rwneg62_10 in62_10 sn62_10 202000.000000
Rwneg63_1 in63_1 sn63_1 202000.000000
Rwneg63_2 in63_2 sn63_2 202000.000000
Rwneg63_3 in63_3 sn63_3 202000.000000
Rwneg63_4 in63_4 sn63_4 78000.000000
Rwneg63_5 in63_5 sn63_5 78000.000000
Rwneg63_6 in63_6 sn63_6 202000.000000
Rwneg63_7 in63_7 sn63_7 202000.000000
Rwneg63_8 in63_8 sn63_8 78000.000000
Rwneg63_9 in63_9 sn63_9 202000.000000
Rwneg63_10 in63_10 sn63_10 202000.000000
Rwneg64_1 in64_1 sn64_1 202000.000000
Rwneg64_2 in64_2 sn64_2 202000.000000
Rwneg64_3 in64_3 sn64_3 202000.000000
Rwneg64_4 in64_4 sn64_4 202000.000000
Rwneg64_5 in64_5 sn64_5 202000.000000
Rwneg64_6 in64_6 sn64_6 202000.000000
Rwneg64_7 in64_7 sn64_7 202000.000000
Rwneg64_8 in64_8 sn64_8 202000.000000
Rwneg64_9 in64_9 sn64_9 202000.000000
Rwneg64_10 in64_10 sn64_10 202000.000000
Rwneg65_1 in65_1 sn65_1 202000.000000
Rwneg65_2 in65_2 sn65_2 202000.000000
Rwneg65_3 in65_3 sn65_3 78000.000000
Rwneg65_4 in65_4 sn65_4 202000.000000
Rwneg65_5 in65_5 sn65_5 202000.000000
Rwneg65_6 in65_6 sn65_6 202000.000000
Rwneg65_7 in65_7 sn65_7 202000.000000
Rwneg65_8 in65_8 sn65_8 78000.000000
Rwneg65_9 in65_9 sn65_9 78000.000000
Rwneg65_10 in65_10 sn65_10 202000.000000
Rwneg66_1 in66_1 sn66_1 78000.000000
Rwneg66_2 in66_2 sn66_2 78000.000000
Rwneg66_3 in66_3 sn66_3 202000.000000
Rwneg66_4 in66_4 sn66_4 78000.000000
Rwneg66_5 in66_5 sn66_5 202000.000000
Rwneg66_6 in66_6 sn66_6 202000.000000
Rwneg66_7 in66_7 sn66_7 202000.000000
Rwneg66_8 in66_8 sn66_8 202000.000000
Rwneg66_9 in66_9 sn66_9 202000.000000
Rwneg66_10 in66_10 sn66_10 78000.000000
Rwneg67_1 in67_1 sn67_1 78000.000000
Rwneg67_2 in67_2 sn67_2 202000.000000
Rwneg67_3 in67_3 sn67_3 202000.000000
Rwneg67_4 in67_4 sn67_4 202000.000000
Rwneg67_5 in67_5 sn67_5 202000.000000
Rwneg67_6 in67_6 sn67_6 78000.000000
Rwneg67_7 in67_7 sn67_7 202000.000000
Rwneg67_8 in67_8 sn67_8 78000.000000
Rwneg67_9 in67_9 sn67_9 202000.000000
Rwneg67_10 in67_10 sn67_10 202000.000000
Rwneg68_1 in68_1 sn68_1 78000.000000
Rwneg68_2 in68_2 sn68_2 78000.000000
Rwneg68_3 in68_3 sn68_3 202000.000000
Rwneg68_4 in68_4 sn68_4 78000.000000
Rwneg68_5 in68_5 sn68_5 202000.000000
Rwneg68_6 in68_6 sn68_6 202000.000000
Rwneg68_7 in68_7 sn68_7 202000.000000
Rwneg68_8 in68_8 sn68_8 78000.000000
Rwneg68_9 in68_9 sn68_9 78000.000000
Rwneg68_10 in68_10 sn68_10 202000.000000
Rwneg69_1 in69_1 sn69_1 202000.000000
Rwneg69_2 in69_2 sn69_2 78000.000000
Rwneg69_3 in69_3 sn69_3 78000.000000
Rwneg69_4 in69_4 sn69_4 78000.000000
Rwneg69_5 in69_5 sn69_5 202000.000000
Rwneg69_6 in69_6 sn69_6 202000.000000
Rwneg69_7 in69_7 sn69_7 78000.000000
Rwneg69_8 in69_8 sn69_8 78000.000000
Rwneg69_9 in69_9 sn69_9 202000.000000
Rwneg69_10 in69_10 sn69_10 202000.000000
Rwneg70_1 in70_1 sn70_1 202000.000000
Rwneg70_2 in70_2 sn70_2 78000.000000
Rwneg70_3 in70_3 sn70_3 78000.000000
Rwneg70_4 in70_4 sn70_4 202000.000000
Rwneg70_5 in70_5 sn70_5 202000.000000
Rwneg70_6 in70_6 sn70_6 202000.000000
Rwneg70_7 in70_7 sn70_7 78000.000000
Rwneg70_8 in70_8 sn70_8 202000.000000
Rwneg70_9 in70_9 sn70_9 202000.000000
Rwneg70_10 in70_10 sn70_10 78000.000000
Rwneg71_1 in71_1 sn71_1 202000.000000
Rwneg71_2 in71_2 sn71_2 202000.000000
Rwneg71_3 in71_3 sn71_3 78000.000000
Rwneg71_4 in71_4 sn71_4 78000.000000
Rwneg71_5 in71_5 sn71_5 78000.000000
Rwneg71_6 in71_6 sn71_6 202000.000000
Rwneg71_7 in71_7 sn71_7 202000.000000
Rwneg71_8 in71_8 sn71_8 78000.000000
Rwneg71_9 in71_9 sn71_9 202000.000000
Rwneg71_10 in71_10 sn71_10 202000.000000
Rwneg72_1 in72_1 sn72_1 202000.000000
Rwneg72_2 in72_2 sn72_2 202000.000000
Rwneg72_3 in72_3 sn72_3 202000.000000
Rwneg72_4 in72_4 sn72_4 202000.000000
Rwneg72_5 in72_5 sn72_5 202000.000000
Rwneg72_6 in72_6 sn72_6 202000.000000
Rwneg72_7 in72_7 sn72_7 78000.000000
Rwneg72_8 in72_8 sn72_8 202000.000000
Rwneg72_9 in72_9 sn72_9 202000.000000
Rwneg72_10 in72_10 sn72_10 202000.000000
Rwneg73_1 in73_1 sn73_1 78000.000000
Rwneg73_2 in73_2 sn73_2 202000.000000
Rwneg73_3 in73_3 sn73_3 78000.000000
Rwneg73_4 in73_4 sn73_4 78000.000000
Rwneg73_5 in73_5 sn73_5 202000.000000
Rwneg73_6 in73_6 sn73_6 202000.000000
Rwneg73_7 in73_7 sn73_7 78000.000000
Rwneg73_8 in73_8 sn73_8 202000.000000
Rwneg73_9 in73_9 sn73_9 202000.000000
Rwneg73_10 in73_10 sn73_10 202000.000000
Rwneg74_1 in74_1 sn74_1 78000.000000
Rwneg74_2 in74_2 sn74_2 202000.000000
Rwneg74_3 in74_3 sn74_3 202000.000000
Rwneg74_4 in74_4 sn74_4 78000.000000
Rwneg74_5 in74_5 sn74_5 202000.000000
Rwneg74_6 in74_6 sn74_6 78000.000000
Rwneg74_7 in74_7 sn74_7 78000.000000
Rwneg74_8 in74_8 sn74_8 202000.000000
Rwneg74_9 in74_9 sn74_9 202000.000000
Rwneg74_10 in74_10 sn74_10 202000.000000
Rwneg75_1 in75_1 sn75_1 202000.000000
Rwneg75_2 in75_2 sn75_2 202000.000000
Rwneg75_3 in75_3 sn75_3 202000.000000
Rwneg75_4 in75_4 sn75_4 202000.000000
Rwneg75_5 in75_5 sn75_5 78000.000000
Rwneg75_6 in75_6 sn75_6 78000.000000
Rwneg75_7 in75_7 sn75_7 78000.000000
Rwneg75_8 in75_8 sn75_8 78000.000000
Rwneg75_9 in75_9 sn75_9 202000.000000
Rwneg75_10 in75_10 sn75_10 202000.000000
Rwneg76_1 in76_1 sn76_1 202000.000000
Rwneg76_2 in76_2 sn76_2 202000.000000
Rwneg76_3 in76_3 sn76_3 202000.000000
Rwneg76_4 in76_4 sn76_4 78000.000000
Rwneg76_5 in76_5 sn76_5 202000.000000
Rwneg76_6 in76_6 sn76_6 78000.000000
Rwneg76_7 in76_7 sn76_7 202000.000000
Rwneg76_8 in76_8 sn76_8 202000.000000
Rwneg76_9 in76_9 sn76_9 202000.000000
Rwneg76_10 in76_10 sn76_10 202000.000000
Rwneg77_1 in77_1 sn77_1 78000.000000
Rwneg77_2 in77_2 sn77_2 202000.000000
Rwneg77_3 in77_3 sn77_3 78000.000000
Rwneg77_4 in77_4 sn77_4 202000.000000
Rwneg77_5 in77_5 sn77_5 78000.000000
Rwneg77_6 in77_6 sn77_6 202000.000000
Rwneg77_7 in77_7 sn77_7 202000.000000
Rwneg77_8 in77_8 sn77_8 78000.000000
Rwneg77_9 in77_9 sn77_9 202000.000000
Rwneg77_10 in77_10 sn77_10 202000.000000
Rwneg78_1 in78_1 sn78_1 78000.000000
Rwneg78_2 in78_2 sn78_2 78000.000000
Rwneg78_3 in78_3 sn78_3 202000.000000
Rwneg78_4 in78_4 sn78_4 78000.000000
Rwneg78_5 in78_5 sn78_5 78000.000000
Rwneg78_6 in78_6 sn78_6 78000.000000
Rwneg78_7 in78_7 sn78_7 78000.000000
Rwneg78_8 in78_8 sn78_8 202000.000000
Rwneg78_9 in78_9 sn78_9 78000.000000
Rwneg78_10 in78_10 sn78_10 78000.000000
Rwneg79_1 in79_1 sn79_1 202000.000000
Rwneg79_2 in79_2 sn79_2 202000.000000
Rwneg79_3 in79_3 sn79_3 78000.000000
Rwneg79_4 in79_4 sn79_4 78000.000000
Rwneg79_5 in79_5 sn79_5 202000.000000
Rwneg79_6 in79_6 sn79_6 202000.000000
Rwneg79_7 in79_7 sn79_7 202000.000000
Rwneg79_8 in79_8 sn79_8 78000.000000
Rwneg79_9 in79_9 sn79_9 202000.000000
Rwneg79_10 in79_10 sn79_10 202000.000000
Rwneg80_1 in80_1 sn80_1 202000.000000
Rwneg80_2 in80_2 sn80_2 78000.000000
Rwneg80_3 in80_3 sn80_3 78000.000000
Rwneg80_4 in80_4 sn80_4 202000.000000
Rwneg80_5 in80_5 sn80_5 78000.000000
Rwneg80_6 in80_6 sn80_6 202000.000000
Rwneg80_7 in80_7 sn80_7 202000.000000
Rwneg80_8 in80_8 sn80_8 202000.000000
Rwneg80_9 in80_9 sn80_9 202000.000000
Rwneg80_10 in80_10 sn80_10 202000.000000
Rwneg81_1 in81_1 sn81_1 202000.000000
Rwneg81_2 in81_2 sn81_2 202000.000000
Rwneg81_3 in81_3 sn81_3 78000.000000
Rwneg81_4 in81_4 sn81_4 202000.000000
Rwneg81_5 in81_5 sn81_5 78000.000000
Rwneg81_6 in81_6 sn81_6 202000.000000
Rwneg81_7 in81_7 sn81_7 202000.000000
Rwneg81_8 in81_8 sn81_8 202000.000000
Rwneg81_9 in81_9 sn81_9 78000.000000
Rwneg81_10 in81_10 sn81_10 202000.000000
Rwneg82_1 in82_1 sn82_1 202000.000000
Rwneg82_2 in82_2 sn82_2 78000.000000
Rwneg82_3 in82_3 sn82_3 202000.000000
Rwneg82_4 in82_4 sn82_4 78000.000000
Rwneg82_5 in82_5 sn82_5 202000.000000
Rwneg82_6 in82_6 sn82_6 202000.000000
Rwneg82_7 in82_7 sn82_7 202000.000000
Rwneg82_8 in82_8 sn82_8 202000.000000
Rwneg82_9 in82_9 sn82_9 202000.000000
Rwneg82_10 in82_10 sn82_10 202000.000000
Rwneg83_1 in83_1 sn83_1 78000.000000
Rwneg83_2 in83_2 sn83_2 202000.000000
Rwneg83_3 in83_3 sn83_3 202000.000000
Rwneg83_4 in83_4 sn83_4 202000.000000
Rwneg83_5 in83_5 sn83_5 78000.000000
Rwneg83_6 in83_6 sn83_6 78000.000000
Rwneg83_7 in83_7 sn83_7 202000.000000
Rwneg83_8 in83_8 sn83_8 202000.000000
Rwneg83_9 in83_9 sn83_9 202000.000000
Rwneg83_10 in83_10 sn83_10 202000.000000
Rwneg84_1 in84_1 sn84_1 78000.000000
Rwneg84_2 in84_2 sn84_2 202000.000000
Rwneg84_3 in84_3 sn84_3 202000.000000
Rwneg84_4 in84_4 sn84_4 202000.000000
Rwneg84_5 in84_5 sn84_5 78000.000000
Rwneg84_6 in84_6 sn84_6 202000.000000
Rwneg84_7 in84_7 sn84_7 202000.000000
Rwneg84_8 in84_8 sn84_8 202000.000000
Rwneg84_9 in84_9 sn84_9 202000.000000
Rwneg84_10 in84_10 sn84_10 202000.000000


**********Positive Biases**********

Rbpos1 vd1 sp85_1 78000.000000
Rbpos2 vd2 sp85_2 202000.000000
Rbpos3 vd3 sp85_3 78000.000000
Rbpos4 vd4 sp85_4 78000.000000
Rbpos5 vd5 sp85_5 78000.000000
Rbpos6 vd6 sp85_6 202000.000000
Rbpos7 vd7 sp85_7 78000.000000
Rbpos8 vd8 sp85_8 78000.000000
Rbpos9 vd9 sp85_9 202000.000000
Rbpos10 vd10 sp85_10 78000.000000


**********Negative Biases**********

Rbneg1 vd1 sn85_1 202000.000000
Rbneg2 vd2 sn85_2 78000.000000
Rbneg3 vd3 sn85_3 202000.000000
Rbneg4 vd4 sn85_4 202000.000000
Rbneg5 vd5 sn85_5 202000.000000
Rbneg6 vd6 sn85_6 78000.000000
Rbneg7 vd7 sn85_7 202000.000000
Rbneg8 vd8 sn85_8 202000.000000
Rbneg9 vd9 sn85_9 78000.000000
Rbneg10 vd10 sn85_10 202000.000000


**********Parasitic Resistances for Vertical Lines**********

Rin1_1 in1 in1_1 9.241569
Rin1_2 in1_1 in1_2 9.241569
Rin1_3 in1_2 in1_3 9.241569
Rin1_4 in1_3 in1_4 9.241569
Rin1_5 in1_4 in1_5 9.241569
Rin1_6 in1_5 in1_6 9.241569
Rin1_7 in1_6 in1_7 9.241569
Rin1_8 in1_7 in1_8 9.241569
Rin1_9 in1_8 in1_9 9.241569
Rin1_10 in1_9 in1_10 9.241569
Rin2_1 in2 in2_1 9.241569
Rin2_2 in2_1 in2_2 9.241569
Rin2_3 in2_2 in2_3 9.241569
Rin2_4 in2_3 in2_4 9.241569
Rin2_5 in2_4 in2_5 9.241569
Rin2_6 in2_5 in2_6 9.241569
Rin2_7 in2_6 in2_7 9.241569
Rin2_8 in2_7 in2_8 9.241569
Rin2_9 in2_8 in2_9 9.241569
Rin2_10 in2_9 in2_10 9.241569
Rin3_1 in3 in3_1 9.241569
Rin3_2 in3_1 in3_2 9.241569
Rin3_3 in3_2 in3_3 9.241569
Rin3_4 in3_3 in3_4 9.241569
Rin3_5 in3_4 in3_5 9.241569
Rin3_6 in3_5 in3_6 9.241569
Rin3_7 in3_6 in3_7 9.241569
Rin3_8 in3_7 in3_8 9.241569
Rin3_9 in3_8 in3_9 9.241569
Rin3_10 in3_9 in3_10 9.241569
Rin4_1 in4 in4_1 9.241569
Rin4_2 in4_1 in4_2 9.241569
Rin4_3 in4_2 in4_3 9.241569
Rin4_4 in4_3 in4_4 9.241569
Rin4_5 in4_4 in4_5 9.241569
Rin4_6 in4_5 in4_6 9.241569
Rin4_7 in4_6 in4_7 9.241569
Rin4_8 in4_7 in4_8 9.241569
Rin4_9 in4_8 in4_9 9.241569
Rin4_10 in4_9 in4_10 9.241569
Rin5_1 in5 in5_1 9.241569
Rin5_2 in5_1 in5_2 9.241569
Rin5_3 in5_2 in5_3 9.241569
Rin5_4 in5_3 in5_4 9.241569
Rin5_5 in5_4 in5_5 9.241569
Rin5_6 in5_5 in5_6 9.241569
Rin5_7 in5_6 in5_7 9.241569
Rin5_8 in5_7 in5_8 9.241569
Rin5_9 in5_8 in5_9 9.241569
Rin5_10 in5_9 in5_10 9.241569
Rin6_1 in6 in6_1 9.241569
Rin6_2 in6_1 in6_2 9.241569
Rin6_3 in6_2 in6_3 9.241569
Rin6_4 in6_3 in6_4 9.241569
Rin6_5 in6_4 in6_5 9.241569
Rin6_6 in6_5 in6_6 9.241569
Rin6_7 in6_6 in6_7 9.241569
Rin6_8 in6_7 in6_8 9.241569
Rin6_9 in6_8 in6_9 9.241569
Rin6_10 in6_9 in6_10 9.241569
Rin7_1 in7 in7_1 9.241569
Rin7_2 in7_1 in7_2 9.241569
Rin7_3 in7_2 in7_3 9.241569
Rin7_4 in7_3 in7_4 9.241569
Rin7_5 in7_4 in7_5 9.241569
Rin7_6 in7_5 in7_6 9.241569
Rin7_7 in7_6 in7_7 9.241569
Rin7_8 in7_7 in7_8 9.241569
Rin7_9 in7_8 in7_9 9.241569
Rin7_10 in7_9 in7_10 9.241569
Rin8_1 in8 in8_1 9.241569
Rin8_2 in8_1 in8_2 9.241569
Rin8_3 in8_2 in8_3 9.241569
Rin8_4 in8_3 in8_4 9.241569
Rin8_5 in8_4 in8_5 9.241569
Rin8_6 in8_5 in8_6 9.241569
Rin8_7 in8_6 in8_7 9.241569
Rin8_8 in8_7 in8_8 9.241569
Rin8_9 in8_8 in8_9 9.241569
Rin8_10 in8_9 in8_10 9.241569
Rin9_1 in9 in9_1 9.241569
Rin9_2 in9_1 in9_2 9.241569
Rin9_3 in9_2 in9_3 9.241569
Rin9_4 in9_3 in9_4 9.241569
Rin9_5 in9_4 in9_5 9.241569
Rin9_6 in9_5 in9_6 9.241569
Rin9_7 in9_6 in9_7 9.241569
Rin9_8 in9_7 in9_8 9.241569
Rin9_9 in9_8 in9_9 9.241569
Rin9_10 in9_9 in9_10 9.241569
Rin10_1 in10 in10_1 9.241569
Rin10_2 in10_1 in10_2 9.241569
Rin10_3 in10_2 in10_3 9.241569
Rin10_4 in10_3 in10_4 9.241569
Rin10_5 in10_4 in10_5 9.241569
Rin10_6 in10_5 in10_6 9.241569
Rin10_7 in10_6 in10_7 9.241569
Rin10_8 in10_7 in10_8 9.241569
Rin10_9 in10_8 in10_9 9.241569
Rin10_10 in10_9 in10_10 9.241569
Rin11_1 in11 in11_1 9.241569
Rin11_2 in11_1 in11_2 9.241569
Rin11_3 in11_2 in11_3 9.241569
Rin11_4 in11_3 in11_4 9.241569
Rin11_5 in11_4 in11_5 9.241569
Rin11_6 in11_5 in11_6 9.241569
Rin11_7 in11_6 in11_7 9.241569
Rin11_8 in11_7 in11_8 9.241569
Rin11_9 in11_8 in11_9 9.241569
Rin11_10 in11_9 in11_10 9.241569
Rin12_1 in12 in12_1 9.241569
Rin12_2 in12_1 in12_2 9.241569
Rin12_3 in12_2 in12_3 9.241569
Rin12_4 in12_3 in12_4 9.241569
Rin12_5 in12_4 in12_5 9.241569
Rin12_6 in12_5 in12_6 9.241569
Rin12_7 in12_6 in12_7 9.241569
Rin12_8 in12_7 in12_8 9.241569
Rin12_9 in12_8 in12_9 9.241569
Rin12_10 in12_9 in12_10 9.241569
Rin13_1 in13 in13_1 9.241569
Rin13_2 in13_1 in13_2 9.241569
Rin13_3 in13_2 in13_3 9.241569
Rin13_4 in13_3 in13_4 9.241569
Rin13_5 in13_4 in13_5 9.241569
Rin13_6 in13_5 in13_6 9.241569
Rin13_7 in13_6 in13_7 9.241569
Rin13_8 in13_7 in13_8 9.241569
Rin13_9 in13_8 in13_9 9.241569
Rin13_10 in13_9 in13_10 9.241569
Rin14_1 in14 in14_1 9.241569
Rin14_2 in14_1 in14_2 9.241569
Rin14_3 in14_2 in14_3 9.241569
Rin14_4 in14_3 in14_4 9.241569
Rin14_5 in14_4 in14_5 9.241569
Rin14_6 in14_5 in14_6 9.241569
Rin14_7 in14_6 in14_7 9.241569
Rin14_8 in14_7 in14_8 9.241569
Rin14_9 in14_8 in14_9 9.241569
Rin14_10 in14_9 in14_10 9.241569
Rin15_1 in15 in15_1 9.241569
Rin15_2 in15_1 in15_2 9.241569
Rin15_3 in15_2 in15_3 9.241569
Rin15_4 in15_3 in15_4 9.241569
Rin15_5 in15_4 in15_5 9.241569
Rin15_6 in15_5 in15_6 9.241569
Rin15_7 in15_6 in15_7 9.241569
Rin15_8 in15_7 in15_8 9.241569
Rin15_9 in15_8 in15_9 9.241569
Rin15_10 in15_9 in15_10 9.241569
Rin16_1 in16 in16_1 9.241569
Rin16_2 in16_1 in16_2 9.241569
Rin16_3 in16_2 in16_3 9.241569
Rin16_4 in16_3 in16_4 9.241569
Rin16_5 in16_4 in16_5 9.241569
Rin16_6 in16_5 in16_6 9.241569
Rin16_7 in16_6 in16_7 9.241569
Rin16_8 in16_7 in16_8 9.241569
Rin16_9 in16_8 in16_9 9.241569
Rin16_10 in16_9 in16_10 9.241569
Rin17_1 in17 in17_1 9.241569
Rin17_2 in17_1 in17_2 9.241569
Rin17_3 in17_2 in17_3 9.241569
Rin17_4 in17_3 in17_4 9.241569
Rin17_5 in17_4 in17_5 9.241569
Rin17_6 in17_5 in17_6 9.241569
Rin17_7 in17_6 in17_7 9.241569
Rin17_8 in17_7 in17_8 9.241569
Rin17_9 in17_8 in17_9 9.241569
Rin17_10 in17_9 in17_10 9.241569
Rin18_1 in18 in18_1 9.241569
Rin18_2 in18_1 in18_2 9.241569
Rin18_3 in18_2 in18_3 9.241569
Rin18_4 in18_3 in18_4 9.241569
Rin18_5 in18_4 in18_5 9.241569
Rin18_6 in18_5 in18_6 9.241569
Rin18_7 in18_6 in18_7 9.241569
Rin18_8 in18_7 in18_8 9.241569
Rin18_9 in18_8 in18_9 9.241569
Rin18_10 in18_9 in18_10 9.241569
Rin19_1 in19 in19_1 9.241569
Rin19_2 in19_1 in19_2 9.241569
Rin19_3 in19_2 in19_3 9.241569
Rin19_4 in19_3 in19_4 9.241569
Rin19_5 in19_4 in19_5 9.241569
Rin19_6 in19_5 in19_6 9.241569
Rin19_7 in19_6 in19_7 9.241569
Rin19_8 in19_7 in19_8 9.241569
Rin19_9 in19_8 in19_9 9.241569
Rin19_10 in19_9 in19_10 9.241569
Rin20_1 in20 in20_1 9.241569
Rin20_2 in20_1 in20_2 9.241569
Rin20_3 in20_2 in20_3 9.241569
Rin20_4 in20_3 in20_4 9.241569
Rin20_5 in20_4 in20_5 9.241569
Rin20_6 in20_5 in20_6 9.241569
Rin20_7 in20_6 in20_7 9.241569
Rin20_8 in20_7 in20_8 9.241569
Rin20_9 in20_8 in20_9 9.241569
Rin20_10 in20_9 in20_10 9.241569
Rin21_1 in21 in21_1 9.241569
Rin21_2 in21_1 in21_2 9.241569
Rin21_3 in21_2 in21_3 9.241569
Rin21_4 in21_3 in21_4 9.241569
Rin21_5 in21_4 in21_5 9.241569
Rin21_6 in21_5 in21_6 9.241569
Rin21_7 in21_6 in21_7 9.241569
Rin21_8 in21_7 in21_8 9.241569
Rin21_9 in21_8 in21_9 9.241569
Rin21_10 in21_9 in21_10 9.241569
Rin22_1 in22 in22_1 9.241569
Rin22_2 in22_1 in22_2 9.241569
Rin22_3 in22_2 in22_3 9.241569
Rin22_4 in22_3 in22_4 9.241569
Rin22_5 in22_4 in22_5 9.241569
Rin22_6 in22_5 in22_6 9.241569
Rin22_7 in22_6 in22_7 9.241569
Rin22_8 in22_7 in22_8 9.241569
Rin22_9 in22_8 in22_9 9.241569
Rin22_10 in22_9 in22_10 9.241569
Rin23_1 in23 in23_1 9.241569
Rin23_2 in23_1 in23_2 9.241569
Rin23_3 in23_2 in23_3 9.241569
Rin23_4 in23_3 in23_4 9.241569
Rin23_5 in23_4 in23_5 9.241569
Rin23_6 in23_5 in23_6 9.241569
Rin23_7 in23_6 in23_7 9.241569
Rin23_8 in23_7 in23_8 9.241569
Rin23_9 in23_8 in23_9 9.241569
Rin23_10 in23_9 in23_10 9.241569
Rin24_1 in24 in24_1 9.241569
Rin24_2 in24_1 in24_2 9.241569
Rin24_3 in24_2 in24_3 9.241569
Rin24_4 in24_3 in24_4 9.241569
Rin24_5 in24_4 in24_5 9.241569
Rin24_6 in24_5 in24_6 9.241569
Rin24_7 in24_6 in24_7 9.241569
Rin24_8 in24_7 in24_8 9.241569
Rin24_9 in24_8 in24_9 9.241569
Rin24_10 in24_9 in24_10 9.241569
Rin25_1 in25 in25_1 9.241569
Rin25_2 in25_1 in25_2 9.241569
Rin25_3 in25_2 in25_3 9.241569
Rin25_4 in25_3 in25_4 9.241569
Rin25_5 in25_4 in25_5 9.241569
Rin25_6 in25_5 in25_6 9.241569
Rin25_7 in25_6 in25_7 9.241569
Rin25_8 in25_7 in25_8 9.241569
Rin25_9 in25_8 in25_9 9.241569
Rin25_10 in25_9 in25_10 9.241569
Rin26_1 in26 in26_1 9.241569
Rin26_2 in26_1 in26_2 9.241569
Rin26_3 in26_2 in26_3 9.241569
Rin26_4 in26_3 in26_4 9.241569
Rin26_5 in26_4 in26_5 9.241569
Rin26_6 in26_5 in26_6 9.241569
Rin26_7 in26_6 in26_7 9.241569
Rin26_8 in26_7 in26_8 9.241569
Rin26_9 in26_8 in26_9 9.241569
Rin26_10 in26_9 in26_10 9.241569
Rin27_1 in27 in27_1 9.241569
Rin27_2 in27_1 in27_2 9.241569
Rin27_3 in27_2 in27_3 9.241569
Rin27_4 in27_3 in27_4 9.241569
Rin27_5 in27_4 in27_5 9.241569
Rin27_6 in27_5 in27_6 9.241569
Rin27_7 in27_6 in27_7 9.241569
Rin27_8 in27_7 in27_8 9.241569
Rin27_9 in27_8 in27_9 9.241569
Rin27_10 in27_9 in27_10 9.241569
Rin28_1 in28 in28_1 9.241569
Rin28_2 in28_1 in28_2 9.241569
Rin28_3 in28_2 in28_3 9.241569
Rin28_4 in28_3 in28_4 9.241569
Rin28_5 in28_4 in28_5 9.241569
Rin28_6 in28_5 in28_6 9.241569
Rin28_7 in28_6 in28_7 9.241569
Rin28_8 in28_7 in28_8 9.241569
Rin28_9 in28_8 in28_9 9.241569
Rin28_10 in28_9 in28_10 9.241569
Rin29_1 in29 in29_1 9.241569
Rin29_2 in29_1 in29_2 9.241569
Rin29_3 in29_2 in29_3 9.241569
Rin29_4 in29_3 in29_4 9.241569
Rin29_5 in29_4 in29_5 9.241569
Rin29_6 in29_5 in29_6 9.241569
Rin29_7 in29_6 in29_7 9.241569
Rin29_8 in29_7 in29_8 9.241569
Rin29_9 in29_8 in29_9 9.241569
Rin29_10 in29_9 in29_10 9.241569
Rin30_1 in30 in30_1 9.241569
Rin30_2 in30_1 in30_2 9.241569
Rin30_3 in30_2 in30_3 9.241569
Rin30_4 in30_3 in30_4 9.241569
Rin30_5 in30_4 in30_5 9.241569
Rin30_6 in30_5 in30_6 9.241569
Rin30_7 in30_6 in30_7 9.241569
Rin30_8 in30_7 in30_8 9.241569
Rin30_9 in30_8 in30_9 9.241569
Rin30_10 in30_9 in30_10 9.241569
Rin31_1 in31 in31_1 9.241569
Rin31_2 in31_1 in31_2 9.241569
Rin31_3 in31_2 in31_3 9.241569
Rin31_4 in31_3 in31_4 9.241569
Rin31_5 in31_4 in31_5 9.241569
Rin31_6 in31_5 in31_6 9.241569
Rin31_7 in31_6 in31_7 9.241569
Rin31_8 in31_7 in31_8 9.241569
Rin31_9 in31_8 in31_9 9.241569
Rin31_10 in31_9 in31_10 9.241569
Rin32_1 in32 in32_1 9.241569
Rin32_2 in32_1 in32_2 9.241569
Rin32_3 in32_2 in32_3 9.241569
Rin32_4 in32_3 in32_4 9.241569
Rin32_5 in32_4 in32_5 9.241569
Rin32_6 in32_5 in32_6 9.241569
Rin32_7 in32_6 in32_7 9.241569
Rin32_8 in32_7 in32_8 9.241569
Rin32_9 in32_8 in32_9 9.241569
Rin32_10 in32_9 in32_10 9.241569
Rin33_1 in33 in33_1 9.241569
Rin33_2 in33_1 in33_2 9.241569
Rin33_3 in33_2 in33_3 9.241569
Rin33_4 in33_3 in33_4 9.241569
Rin33_5 in33_4 in33_5 9.241569
Rin33_6 in33_5 in33_6 9.241569
Rin33_7 in33_6 in33_7 9.241569
Rin33_8 in33_7 in33_8 9.241569
Rin33_9 in33_8 in33_9 9.241569
Rin33_10 in33_9 in33_10 9.241569
Rin34_1 in34 in34_1 9.241569
Rin34_2 in34_1 in34_2 9.241569
Rin34_3 in34_2 in34_3 9.241569
Rin34_4 in34_3 in34_4 9.241569
Rin34_5 in34_4 in34_5 9.241569
Rin34_6 in34_5 in34_6 9.241569
Rin34_7 in34_6 in34_7 9.241569
Rin34_8 in34_7 in34_8 9.241569
Rin34_9 in34_8 in34_9 9.241569
Rin34_10 in34_9 in34_10 9.241569
Rin35_1 in35 in35_1 9.241569
Rin35_2 in35_1 in35_2 9.241569
Rin35_3 in35_2 in35_3 9.241569
Rin35_4 in35_3 in35_4 9.241569
Rin35_5 in35_4 in35_5 9.241569
Rin35_6 in35_5 in35_6 9.241569
Rin35_7 in35_6 in35_7 9.241569
Rin35_8 in35_7 in35_8 9.241569
Rin35_9 in35_8 in35_9 9.241569
Rin35_10 in35_9 in35_10 9.241569
Rin36_1 in36 in36_1 9.241569
Rin36_2 in36_1 in36_2 9.241569
Rin36_3 in36_2 in36_3 9.241569
Rin36_4 in36_3 in36_4 9.241569
Rin36_5 in36_4 in36_5 9.241569
Rin36_6 in36_5 in36_6 9.241569
Rin36_7 in36_6 in36_7 9.241569
Rin36_8 in36_7 in36_8 9.241569
Rin36_9 in36_8 in36_9 9.241569
Rin36_10 in36_9 in36_10 9.241569
Rin37_1 in37 in37_1 9.241569
Rin37_2 in37_1 in37_2 9.241569
Rin37_3 in37_2 in37_3 9.241569
Rin37_4 in37_3 in37_4 9.241569
Rin37_5 in37_4 in37_5 9.241569
Rin37_6 in37_5 in37_6 9.241569
Rin37_7 in37_6 in37_7 9.241569
Rin37_8 in37_7 in37_8 9.241569
Rin37_9 in37_8 in37_9 9.241569
Rin37_10 in37_9 in37_10 9.241569
Rin38_1 in38 in38_1 9.241569
Rin38_2 in38_1 in38_2 9.241569
Rin38_3 in38_2 in38_3 9.241569
Rin38_4 in38_3 in38_4 9.241569
Rin38_5 in38_4 in38_5 9.241569
Rin38_6 in38_5 in38_6 9.241569
Rin38_7 in38_6 in38_7 9.241569
Rin38_8 in38_7 in38_8 9.241569
Rin38_9 in38_8 in38_9 9.241569
Rin38_10 in38_9 in38_10 9.241569
Rin39_1 in39 in39_1 9.241569
Rin39_2 in39_1 in39_2 9.241569
Rin39_3 in39_2 in39_3 9.241569
Rin39_4 in39_3 in39_4 9.241569
Rin39_5 in39_4 in39_5 9.241569
Rin39_6 in39_5 in39_6 9.241569
Rin39_7 in39_6 in39_7 9.241569
Rin39_8 in39_7 in39_8 9.241569
Rin39_9 in39_8 in39_9 9.241569
Rin39_10 in39_9 in39_10 9.241569
Rin40_1 in40 in40_1 9.241569
Rin40_2 in40_1 in40_2 9.241569
Rin40_3 in40_2 in40_3 9.241569
Rin40_4 in40_3 in40_4 9.241569
Rin40_5 in40_4 in40_5 9.241569
Rin40_6 in40_5 in40_6 9.241569
Rin40_7 in40_6 in40_7 9.241569
Rin40_8 in40_7 in40_8 9.241569
Rin40_9 in40_8 in40_9 9.241569
Rin40_10 in40_9 in40_10 9.241569
Rin41_1 in41 in41_1 9.241569
Rin41_2 in41_1 in41_2 9.241569
Rin41_3 in41_2 in41_3 9.241569
Rin41_4 in41_3 in41_4 9.241569
Rin41_5 in41_4 in41_5 9.241569
Rin41_6 in41_5 in41_6 9.241569
Rin41_7 in41_6 in41_7 9.241569
Rin41_8 in41_7 in41_8 9.241569
Rin41_9 in41_8 in41_9 9.241569
Rin41_10 in41_9 in41_10 9.241569
Rin42_1 in42 in42_1 9.241569
Rin42_2 in42_1 in42_2 9.241569
Rin42_3 in42_2 in42_3 9.241569
Rin42_4 in42_3 in42_4 9.241569
Rin42_5 in42_4 in42_5 9.241569
Rin42_6 in42_5 in42_6 9.241569
Rin42_7 in42_6 in42_7 9.241569
Rin42_8 in42_7 in42_8 9.241569
Rin42_9 in42_8 in42_9 9.241569
Rin42_10 in42_9 in42_10 9.241569
Rin43_1 in43 in43_1 9.241569
Rin43_2 in43_1 in43_2 9.241569
Rin43_3 in43_2 in43_3 9.241569
Rin43_4 in43_3 in43_4 9.241569
Rin43_5 in43_4 in43_5 9.241569
Rin43_6 in43_5 in43_6 9.241569
Rin43_7 in43_6 in43_7 9.241569
Rin43_8 in43_7 in43_8 9.241569
Rin43_9 in43_8 in43_9 9.241569
Rin43_10 in43_9 in43_10 9.241569
Rin44_1 in44 in44_1 9.241569
Rin44_2 in44_1 in44_2 9.241569
Rin44_3 in44_2 in44_3 9.241569
Rin44_4 in44_3 in44_4 9.241569
Rin44_5 in44_4 in44_5 9.241569
Rin44_6 in44_5 in44_6 9.241569
Rin44_7 in44_6 in44_7 9.241569
Rin44_8 in44_7 in44_8 9.241569
Rin44_9 in44_8 in44_9 9.241569
Rin44_10 in44_9 in44_10 9.241569
Rin45_1 in45 in45_1 9.241569
Rin45_2 in45_1 in45_2 9.241569
Rin45_3 in45_2 in45_3 9.241569
Rin45_4 in45_3 in45_4 9.241569
Rin45_5 in45_4 in45_5 9.241569
Rin45_6 in45_5 in45_6 9.241569
Rin45_7 in45_6 in45_7 9.241569
Rin45_8 in45_7 in45_8 9.241569
Rin45_9 in45_8 in45_9 9.241569
Rin45_10 in45_9 in45_10 9.241569
Rin46_1 in46 in46_1 9.241569
Rin46_2 in46_1 in46_2 9.241569
Rin46_3 in46_2 in46_3 9.241569
Rin46_4 in46_3 in46_4 9.241569
Rin46_5 in46_4 in46_5 9.241569
Rin46_6 in46_5 in46_6 9.241569
Rin46_7 in46_6 in46_7 9.241569
Rin46_8 in46_7 in46_8 9.241569
Rin46_9 in46_8 in46_9 9.241569
Rin46_10 in46_9 in46_10 9.241569
Rin47_1 in47 in47_1 9.241569
Rin47_2 in47_1 in47_2 9.241569
Rin47_3 in47_2 in47_3 9.241569
Rin47_4 in47_3 in47_4 9.241569
Rin47_5 in47_4 in47_5 9.241569
Rin47_6 in47_5 in47_6 9.241569
Rin47_7 in47_6 in47_7 9.241569
Rin47_8 in47_7 in47_8 9.241569
Rin47_9 in47_8 in47_9 9.241569
Rin47_10 in47_9 in47_10 9.241569
Rin48_1 in48 in48_1 9.241569
Rin48_2 in48_1 in48_2 9.241569
Rin48_3 in48_2 in48_3 9.241569
Rin48_4 in48_3 in48_4 9.241569
Rin48_5 in48_4 in48_5 9.241569
Rin48_6 in48_5 in48_6 9.241569
Rin48_7 in48_6 in48_7 9.241569
Rin48_8 in48_7 in48_8 9.241569
Rin48_9 in48_8 in48_9 9.241569
Rin48_10 in48_9 in48_10 9.241569
Rin49_1 in49 in49_1 9.241569
Rin49_2 in49_1 in49_2 9.241569
Rin49_3 in49_2 in49_3 9.241569
Rin49_4 in49_3 in49_4 9.241569
Rin49_5 in49_4 in49_5 9.241569
Rin49_6 in49_5 in49_6 9.241569
Rin49_7 in49_6 in49_7 9.241569
Rin49_8 in49_7 in49_8 9.241569
Rin49_9 in49_8 in49_9 9.241569
Rin49_10 in49_9 in49_10 9.241569
Rin50_1 in50 in50_1 9.241569
Rin50_2 in50_1 in50_2 9.241569
Rin50_3 in50_2 in50_3 9.241569
Rin50_4 in50_3 in50_4 9.241569
Rin50_5 in50_4 in50_5 9.241569
Rin50_6 in50_5 in50_6 9.241569
Rin50_7 in50_6 in50_7 9.241569
Rin50_8 in50_7 in50_8 9.241569
Rin50_9 in50_8 in50_9 9.241569
Rin50_10 in50_9 in50_10 9.241569
Rin51_1 in51 in51_1 9.241569
Rin51_2 in51_1 in51_2 9.241569
Rin51_3 in51_2 in51_3 9.241569
Rin51_4 in51_3 in51_4 9.241569
Rin51_5 in51_4 in51_5 9.241569
Rin51_6 in51_5 in51_6 9.241569
Rin51_7 in51_6 in51_7 9.241569
Rin51_8 in51_7 in51_8 9.241569
Rin51_9 in51_8 in51_9 9.241569
Rin51_10 in51_9 in51_10 9.241569
Rin52_1 in52 in52_1 9.241569
Rin52_2 in52_1 in52_2 9.241569
Rin52_3 in52_2 in52_3 9.241569
Rin52_4 in52_3 in52_4 9.241569
Rin52_5 in52_4 in52_5 9.241569
Rin52_6 in52_5 in52_6 9.241569
Rin52_7 in52_6 in52_7 9.241569
Rin52_8 in52_7 in52_8 9.241569
Rin52_9 in52_8 in52_9 9.241569
Rin52_10 in52_9 in52_10 9.241569
Rin53_1 in53 in53_1 9.241569
Rin53_2 in53_1 in53_2 9.241569
Rin53_3 in53_2 in53_3 9.241569
Rin53_4 in53_3 in53_4 9.241569
Rin53_5 in53_4 in53_5 9.241569
Rin53_6 in53_5 in53_6 9.241569
Rin53_7 in53_6 in53_7 9.241569
Rin53_8 in53_7 in53_8 9.241569
Rin53_9 in53_8 in53_9 9.241569
Rin53_10 in53_9 in53_10 9.241569
Rin54_1 in54 in54_1 9.241569
Rin54_2 in54_1 in54_2 9.241569
Rin54_3 in54_2 in54_3 9.241569
Rin54_4 in54_3 in54_4 9.241569
Rin54_5 in54_4 in54_5 9.241569
Rin54_6 in54_5 in54_6 9.241569
Rin54_7 in54_6 in54_7 9.241569
Rin54_8 in54_7 in54_8 9.241569
Rin54_9 in54_8 in54_9 9.241569
Rin54_10 in54_9 in54_10 9.241569
Rin55_1 in55 in55_1 9.241569
Rin55_2 in55_1 in55_2 9.241569
Rin55_3 in55_2 in55_3 9.241569
Rin55_4 in55_3 in55_4 9.241569
Rin55_5 in55_4 in55_5 9.241569
Rin55_6 in55_5 in55_6 9.241569
Rin55_7 in55_6 in55_7 9.241569
Rin55_8 in55_7 in55_8 9.241569
Rin55_9 in55_8 in55_9 9.241569
Rin55_10 in55_9 in55_10 9.241569
Rin56_1 in56 in56_1 9.241569
Rin56_2 in56_1 in56_2 9.241569
Rin56_3 in56_2 in56_3 9.241569
Rin56_4 in56_3 in56_4 9.241569
Rin56_5 in56_4 in56_5 9.241569
Rin56_6 in56_5 in56_6 9.241569
Rin56_7 in56_6 in56_7 9.241569
Rin56_8 in56_7 in56_8 9.241569
Rin56_9 in56_8 in56_9 9.241569
Rin56_10 in56_9 in56_10 9.241569
Rin57_1 in57 in57_1 9.241569
Rin57_2 in57_1 in57_2 9.241569
Rin57_3 in57_2 in57_3 9.241569
Rin57_4 in57_3 in57_4 9.241569
Rin57_5 in57_4 in57_5 9.241569
Rin57_6 in57_5 in57_6 9.241569
Rin57_7 in57_6 in57_7 9.241569
Rin57_8 in57_7 in57_8 9.241569
Rin57_9 in57_8 in57_9 9.241569
Rin57_10 in57_9 in57_10 9.241569
Rin58_1 in58 in58_1 9.241569
Rin58_2 in58_1 in58_2 9.241569
Rin58_3 in58_2 in58_3 9.241569
Rin58_4 in58_3 in58_4 9.241569
Rin58_5 in58_4 in58_5 9.241569
Rin58_6 in58_5 in58_6 9.241569
Rin58_7 in58_6 in58_7 9.241569
Rin58_8 in58_7 in58_8 9.241569
Rin58_9 in58_8 in58_9 9.241569
Rin58_10 in58_9 in58_10 9.241569
Rin59_1 in59 in59_1 9.241569
Rin59_2 in59_1 in59_2 9.241569
Rin59_3 in59_2 in59_3 9.241569
Rin59_4 in59_3 in59_4 9.241569
Rin59_5 in59_4 in59_5 9.241569
Rin59_6 in59_5 in59_6 9.241569
Rin59_7 in59_6 in59_7 9.241569
Rin59_8 in59_7 in59_8 9.241569
Rin59_9 in59_8 in59_9 9.241569
Rin59_10 in59_9 in59_10 9.241569
Rin60_1 in60 in60_1 9.241569
Rin60_2 in60_1 in60_2 9.241569
Rin60_3 in60_2 in60_3 9.241569
Rin60_4 in60_3 in60_4 9.241569
Rin60_5 in60_4 in60_5 9.241569
Rin60_6 in60_5 in60_6 9.241569
Rin60_7 in60_6 in60_7 9.241569
Rin60_8 in60_7 in60_8 9.241569
Rin60_9 in60_8 in60_9 9.241569
Rin60_10 in60_9 in60_10 9.241569
Rin61_1 in61 in61_1 9.241569
Rin61_2 in61_1 in61_2 9.241569
Rin61_3 in61_2 in61_3 9.241569
Rin61_4 in61_3 in61_4 9.241569
Rin61_5 in61_4 in61_5 9.241569
Rin61_6 in61_5 in61_6 9.241569
Rin61_7 in61_6 in61_7 9.241569
Rin61_8 in61_7 in61_8 9.241569
Rin61_9 in61_8 in61_9 9.241569
Rin61_10 in61_9 in61_10 9.241569
Rin62_1 in62 in62_1 9.241569
Rin62_2 in62_1 in62_2 9.241569
Rin62_3 in62_2 in62_3 9.241569
Rin62_4 in62_3 in62_4 9.241569
Rin62_5 in62_4 in62_5 9.241569
Rin62_6 in62_5 in62_6 9.241569
Rin62_7 in62_6 in62_7 9.241569
Rin62_8 in62_7 in62_8 9.241569
Rin62_9 in62_8 in62_9 9.241569
Rin62_10 in62_9 in62_10 9.241569
Rin63_1 in63 in63_1 9.241569
Rin63_2 in63_1 in63_2 9.241569
Rin63_3 in63_2 in63_3 9.241569
Rin63_4 in63_3 in63_4 9.241569
Rin63_5 in63_4 in63_5 9.241569
Rin63_6 in63_5 in63_6 9.241569
Rin63_7 in63_6 in63_7 9.241569
Rin63_8 in63_7 in63_8 9.241569
Rin63_9 in63_8 in63_9 9.241569
Rin63_10 in63_9 in63_10 9.241569
Rin64_1 in64 in64_1 9.241569
Rin64_2 in64_1 in64_2 9.241569
Rin64_3 in64_2 in64_3 9.241569
Rin64_4 in64_3 in64_4 9.241569
Rin64_5 in64_4 in64_5 9.241569
Rin64_6 in64_5 in64_6 9.241569
Rin64_7 in64_6 in64_7 9.241569
Rin64_8 in64_7 in64_8 9.241569
Rin64_9 in64_8 in64_9 9.241569
Rin64_10 in64_9 in64_10 9.241569
Rin65_1 in65 in65_1 9.241569
Rin65_2 in65_1 in65_2 9.241569
Rin65_3 in65_2 in65_3 9.241569
Rin65_4 in65_3 in65_4 9.241569
Rin65_5 in65_4 in65_5 9.241569
Rin65_6 in65_5 in65_6 9.241569
Rin65_7 in65_6 in65_7 9.241569
Rin65_8 in65_7 in65_8 9.241569
Rin65_9 in65_8 in65_9 9.241569
Rin65_10 in65_9 in65_10 9.241569
Rin66_1 in66 in66_1 9.241569
Rin66_2 in66_1 in66_2 9.241569
Rin66_3 in66_2 in66_3 9.241569
Rin66_4 in66_3 in66_4 9.241569
Rin66_5 in66_4 in66_5 9.241569
Rin66_6 in66_5 in66_6 9.241569
Rin66_7 in66_6 in66_7 9.241569
Rin66_8 in66_7 in66_8 9.241569
Rin66_9 in66_8 in66_9 9.241569
Rin66_10 in66_9 in66_10 9.241569
Rin67_1 in67 in67_1 9.241569
Rin67_2 in67_1 in67_2 9.241569
Rin67_3 in67_2 in67_3 9.241569
Rin67_4 in67_3 in67_4 9.241569
Rin67_5 in67_4 in67_5 9.241569
Rin67_6 in67_5 in67_6 9.241569
Rin67_7 in67_6 in67_7 9.241569
Rin67_8 in67_7 in67_8 9.241569
Rin67_9 in67_8 in67_9 9.241569
Rin67_10 in67_9 in67_10 9.241569
Rin68_1 in68 in68_1 9.241569
Rin68_2 in68_1 in68_2 9.241569
Rin68_3 in68_2 in68_3 9.241569
Rin68_4 in68_3 in68_4 9.241569
Rin68_5 in68_4 in68_5 9.241569
Rin68_6 in68_5 in68_6 9.241569
Rin68_7 in68_6 in68_7 9.241569
Rin68_8 in68_7 in68_8 9.241569
Rin68_9 in68_8 in68_9 9.241569
Rin68_10 in68_9 in68_10 9.241569
Rin69_1 in69 in69_1 9.241569
Rin69_2 in69_1 in69_2 9.241569
Rin69_3 in69_2 in69_3 9.241569
Rin69_4 in69_3 in69_4 9.241569
Rin69_5 in69_4 in69_5 9.241569
Rin69_6 in69_5 in69_6 9.241569
Rin69_7 in69_6 in69_7 9.241569
Rin69_8 in69_7 in69_8 9.241569
Rin69_9 in69_8 in69_9 9.241569
Rin69_10 in69_9 in69_10 9.241569
Rin70_1 in70 in70_1 9.241569
Rin70_2 in70_1 in70_2 9.241569
Rin70_3 in70_2 in70_3 9.241569
Rin70_4 in70_3 in70_4 9.241569
Rin70_5 in70_4 in70_5 9.241569
Rin70_6 in70_5 in70_6 9.241569
Rin70_7 in70_6 in70_7 9.241569
Rin70_8 in70_7 in70_8 9.241569
Rin70_9 in70_8 in70_9 9.241569
Rin70_10 in70_9 in70_10 9.241569
Rin71_1 in71 in71_1 9.241569
Rin71_2 in71_1 in71_2 9.241569
Rin71_3 in71_2 in71_3 9.241569
Rin71_4 in71_3 in71_4 9.241569
Rin71_5 in71_4 in71_5 9.241569
Rin71_6 in71_5 in71_6 9.241569
Rin71_7 in71_6 in71_7 9.241569
Rin71_8 in71_7 in71_8 9.241569
Rin71_9 in71_8 in71_9 9.241569
Rin71_10 in71_9 in71_10 9.241569
Rin72_1 in72 in72_1 9.241569
Rin72_2 in72_1 in72_2 9.241569
Rin72_3 in72_2 in72_3 9.241569
Rin72_4 in72_3 in72_4 9.241569
Rin72_5 in72_4 in72_5 9.241569
Rin72_6 in72_5 in72_6 9.241569
Rin72_7 in72_6 in72_7 9.241569
Rin72_8 in72_7 in72_8 9.241569
Rin72_9 in72_8 in72_9 9.241569
Rin72_10 in72_9 in72_10 9.241569
Rin73_1 in73 in73_1 9.241569
Rin73_2 in73_1 in73_2 9.241569
Rin73_3 in73_2 in73_3 9.241569
Rin73_4 in73_3 in73_4 9.241569
Rin73_5 in73_4 in73_5 9.241569
Rin73_6 in73_5 in73_6 9.241569
Rin73_7 in73_6 in73_7 9.241569
Rin73_8 in73_7 in73_8 9.241569
Rin73_9 in73_8 in73_9 9.241569
Rin73_10 in73_9 in73_10 9.241569
Rin74_1 in74 in74_1 9.241569
Rin74_2 in74_1 in74_2 9.241569
Rin74_3 in74_2 in74_3 9.241569
Rin74_4 in74_3 in74_4 9.241569
Rin74_5 in74_4 in74_5 9.241569
Rin74_6 in74_5 in74_6 9.241569
Rin74_7 in74_6 in74_7 9.241569
Rin74_8 in74_7 in74_8 9.241569
Rin74_9 in74_8 in74_9 9.241569
Rin74_10 in74_9 in74_10 9.241569
Rin75_1 in75 in75_1 9.241569
Rin75_2 in75_1 in75_2 9.241569
Rin75_3 in75_2 in75_3 9.241569
Rin75_4 in75_3 in75_4 9.241569
Rin75_5 in75_4 in75_5 9.241569
Rin75_6 in75_5 in75_6 9.241569
Rin75_7 in75_6 in75_7 9.241569
Rin75_8 in75_7 in75_8 9.241569
Rin75_9 in75_8 in75_9 9.241569
Rin75_10 in75_9 in75_10 9.241569
Rin76_1 in76 in76_1 9.241569
Rin76_2 in76_1 in76_2 9.241569
Rin76_3 in76_2 in76_3 9.241569
Rin76_4 in76_3 in76_4 9.241569
Rin76_5 in76_4 in76_5 9.241569
Rin76_6 in76_5 in76_6 9.241569
Rin76_7 in76_6 in76_7 9.241569
Rin76_8 in76_7 in76_8 9.241569
Rin76_9 in76_8 in76_9 9.241569
Rin76_10 in76_9 in76_10 9.241569
Rin77_1 in77 in77_1 9.241569
Rin77_2 in77_1 in77_2 9.241569
Rin77_3 in77_2 in77_3 9.241569
Rin77_4 in77_3 in77_4 9.241569
Rin77_5 in77_4 in77_5 9.241569
Rin77_6 in77_5 in77_6 9.241569
Rin77_7 in77_6 in77_7 9.241569
Rin77_8 in77_7 in77_8 9.241569
Rin77_9 in77_8 in77_9 9.241569
Rin77_10 in77_9 in77_10 9.241569
Rin78_1 in78 in78_1 9.241569
Rin78_2 in78_1 in78_2 9.241569
Rin78_3 in78_2 in78_3 9.241569
Rin78_4 in78_3 in78_4 9.241569
Rin78_5 in78_4 in78_5 9.241569
Rin78_6 in78_5 in78_6 9.241569
Rin78_7 in78_6 in78_7 9.241569
Rin78_8 in78_7 in78_8 9.241569
Rin78_9 in78_8 in78_9 9.241569
Rin78_10 in78_9 in78_10 9.241569
Rin79_1 in79 in79_1 9.241569
Rin79_2 in79_1 in79_2 9.241569
Rin79_3 in79_2 in79_3 9.241569
Rin79_4 in79_3 in79_4 9.241569
Rin79_5 in79_4 in79_5 9.241569
Rin79_6 in79_5 in79_6 9.241569
Rin79_7 in79_6 in79_7 9.241569
Rin79_8 in79_7 in79_8 9.241569
Rin79_9 in79_8 in79_9 9.241569
Rin79_10 in79_9 in79_10 9.241569
Rin80_1 in80 in80_1 9.241569
Rin80_2 in80_1 in80_2 9.241569
Rin80_3 in80_2 in80_3 9.241569
Rin80_4 in80_3 in80_4 9.241569
Rin80_5 in80_4 in80_5 9.241569
Rin80_6 in80_5 in80_6 9.241569
Rin80_7 in80_6 in80_7 9.241569
Rin80_8 in80_7 in80_8 9.241569
Rin80_9 in80_8 in80_9 9.241569
Rin80_10 in80_9 in80_10 9.241569
Rin81_1 in81 in81_1 9.241569
Rin81_2 in81_1 in81_2 9.241569
Rin81_3 in81_2 in81_3 9.241569
Rin81_4 in81_3 in81_4 9.241569
Rin81_5 in81_4 in81_5 9.241569
Rin81_6 in81_5 in81_6 9.241569
Rin81_7 in81_6 in81_7 9.241569
Rin81_8 in81_7 in81_8 9.241569
Rin81_9 in81_8 in81_9 9.241569
Rin81_10 in81_9 in81_10 9.241569
Rin82_1 in82 in82_1 9.241569
Rin82_2 in82_1 in82_2 9.241569
Rin82_3 in82_2 in82_3 9.241569
Rin82_4 in82_3 in82_4 9.241569
Rin82_5 in82_4 in82_5 9.241569
Rin82_6 in82_5 in82_6 9.241569
Rin82_7 in82_6 in82_7 9.241569
Rin82_8 in82_7 in82_8 9.241569
Rin82_9 in82_8 in82_9 9.241569
Rin82_10 in82_9 in82_10 9.241569
Rin83_1 in83 in83_1 9.241569
Rin83_2 in83_1 in83_2 9.241569
Rin83_3 in83_2 in83_3 9.241569
Rin83_4 in83_3 in83_4 9.241569
Rin83_5 in83_4 in83_5 9.241569
Rin83_6 in83_5 in83_6 9.241569
Rin83_7 in83_6 in83_7 9.241569
Rin83_8 in83_7 in83_8 9.241569
Rin83_9 in83_8 in83_9 9.241569
Rin83_10 in83_9 in83_10 9.241569
Rin84_1 in84 in84_1 9.241569
Rin84_2 in84_1 in84_2 9.241569
Rin84_3 in84_2 in84_3 9.241569
Rin84_4 in84_3 in84_4 9.241569
Rin84_5 in84_4 in84_5 9.241569
Rin84_6 in84_5 in84_6 9.241569
Rin84_7 in84_6 in84_7 9.241569
Rin84_8 in84_7 in84_8 9.241569
Rin84_9 in84_8 in84_9 9.241569
Rin84_10 in84_9 in84_10 9.241569
Rbias1 vdd vd1 9.241569
Rbias2 vd1 vd2 9.241569
Rbias3 vd2 vd3 9.241569
Rbias4 vd3 vd4 9.241569
Rbias5 vd4 vd5 9.241569
Rbias6 vd5 vd6 9.241569
Rbias7 vd6 vd7 9.241569
Rbias8 vd7 vd8 9.241569
Rbias9 vd8 vd9 9.241569
Rbias10 vd9 vd10 9.241569


**********Parasitic Resistances for I+ and I- Lines****************

Rsp1_1 sp1_1 sp2_1 11.551961
Rsn1_1 sn1_1 sn2_1 11.551961
Rsp1_2 sp1_2 sp2_2 11.551961
Rsn1_2 sn1_2 sn2_2 11.551961
Rsp1_3 sp1_3 sp2_3 11.551961
Rsn1_3 sn1_3 sn2_3 11.551961
Rsp1_4 sp1_4 sp2_4 11.551961
Rsn1_4 sn1_4 sn2_4 11.551961
Rsp1_5 sp1_5 sp2_5 11.551961
Rsn1_5 sn1_5 sn2_5 11.551961
Rsp1_6 sp1_6 sp2_6 11.551961
Rsn1_6 sn1_6 sn2_6 11.551961
Rsp1_7 sp1_7 sp2_7 11.551961
Rsn1_7 sn1_7 sn2_7 11.551961
Rsp1_8 sp1_8 sp2_8 11.551961
Rsn1_8 sn1_8 sn2_8 11.551961
Rsp1_9 sp1_9 sp2_9 11.551961
Rsn1_9 sn1_9 sn2_9 11.551961
Rsp1_10 sp1_10 sp2_10 11.551961
Rsn1_10 sn1_10 sn2_10 11.551961
Rsp2_1 sp2_1 sp3_1 11.551961
Rsn2_1 sn2_1 sn3_1 11.551961
Rsp2_2 sp2_2 sp3_2 11.551961
Rsn2_2 sn2_2 sn3_2 11.551961
Rsp2_3 sp2_3 sp3_3 11.551961
Rsn2_3 sn2_3 sn3_3 11.551961
Rsp2_4 sp2_4 sp3_4 11.551961
Rsn2_4 sn2_4 sn3_4 11.551961
Rsp2_5 sp2_5 sp3_5 11.551961
Rsn2_5 sn2_5 sn3_5 11.551961
Rsp2_6 sp2_6 sp3_6 11.551961
Rsn2_6 sn2_6 sn3_6 11.551961
Rsp2_7 sp2_7 sp3_7 11.551961
Rsn2_7 sn2_7 sn3_7 11.551961
Rsp2_8 sp2_8 sp3_8 11.551961
Rsn2_8 sn2_8 sn3_8 11.551961
Rsp2_9 sp2_9 sp3_9 11.551961
Rsn2_9 sn2_9 sn3_9 11.551961
Rsp2_10 sp2_10 sp3_10 11.551961
Rsn2_10 sn2_10 sn3_10 11.551961
Rsp3_1 sp3_1 sp4_1 11.551961
Rsn3_1 sn3_1 sn4_1 11.551961
Rsp3_2 sp3_2 sp4_2 11.551961
Rsn3_2 sn3_2 sn4_2 11.551961
Rsp3_3 sp3_3 sp4_3 11.551961
Rsn3_3 sn3_3 sn4_3 11.551961
Rsp3_4 sp3_4 sp4_4 11.551961
Rsn3_4 sn3_4 sn4_4 11.551961
Rsp3_5 sp3_5 sp4_5 11.551961
Rsn3_5 sn3_5 sn4_5 11.551961
Rsp3_6 sp3_6 sp4_6 11.551961
Rsn3_6 sn3_6 sn4_6 11.551961
Rsp3_7 sp3_7 sp4_7 11.551961
Rsn3_7 sn3_7 sn4_7 11.551961
Rsp3_8 sp3_8 sp4_8 11.551961
Rsn3_8 sn3_8 sn4_8 11.551961
Rsp3_9 sp3_9 sp4_9 11.551961
Rsn3_9 sn3_9 sn4_9 11.551961
Rsp3_10 sp3_10 sp4_10 11.551961
Rsn3_10 sn3_10 sn4_10 11.551961
Rsp4_1 sp4_1 sp5_1 11.551961
Rsn4_1 sn4_1 sn5_1 11.551961
Rsp4_2 sp4_2 sp5_2 11.551961
Rsn4_2 sn4_2 sn5_2 11.551961
Rsp4_3 sp4_3 sp5_3 11.551961
Rsn4_3 sn4_3 sn5_3 11.551961
Rsp4_4 sp4_4 sp5_4 11.551961
Rsn4_4 sn4_4 sn5_4 11.551961
Rsp4_5 sp4_5 sp5_5 11.551961
Rsn4_5 sn4_5 sn5_5 11.551961
Rsp4_6 sp4_6 sp5_6 11.551961
Rsn4_6 sn4_6 sn5_6 11.551961
Rsp4_7 sp4_7 sp5_7 11.551961
Rsn4_7 sn4_7 sn5_7 11.551961
Rsp4_8 sp4_8 sp5_8 11.551961
Rsn4_8 sn4_8 sn5_8 11.551961
Rsp4_9 sp4_9 sp5_9 11.551961
Rsn4_9 sn4_9 sn5_9 11.551961
Rsp4_10 sp4_10 sp5_10 11.551961
Rsn4_10 sn4_10 sn5_10 11.551961
Rsp5_1 sp5_1 sp6_1 11.551961
Rsn5_1 sn5_1 sn6_1 11.551961
Rsp5_2 sp5_2 sp6_2 11.551961
Rsn5_2 sn5_2 sn6_2 11.551961
Rsp5_3 sp5_3 sp6_3 11.551961
Rsn5_3 sn5_3 sn6_3 11.551961
Rsp5_4 sp5_4 sp6_4 11.551961
Rsn5_4 sn5_4 sn6_4 11.551961
Rsp5_5 sp5_5 sp6_5 11.551961
Rsn5_5 sn5_5 sn6_5 11.551961
Rsp5_6 sp5_6 sp6_6 11.551961
Rsn5_6 sn5_6 sn6_6 11.551961
Rsp5_7 sp5_7 sp6_7 11.551961
Rsn5_7 sn5_7 sn6_7 11.551961
Rsp5_8 sp5_8 sp6_8 11.551961
Rsn5_8 sn5_8 sn6_8 11.551961
Rsp5_9 sp5_9 sp6_9 11.551961
Rsn5_9 sn5_9 sn6_9 11.551961
Rsp5_10 sp5_10 sp6_10 11.551961
Rsn5_10 sn5_10 sn6_10 11.551961
Rsp6_1 sp6_1 sp7_1 11.551961
Rsn6_1 sn6_1 sn7_1 11.551961
Rsp6_2 sp6_2 sp7_2 11.551961
Rsn6_2 sn6_2 sn7_2 11.551961
Rsp6_3 sp6_3 sp7_3 11.551961
Rsn6_3 sn6_3 sn7_3 11.551961
Rsp6_4 sp6_4 sp7_4 11.551961
Rsn6_4 sn6_4 sn7_4 11.551961
Rsp6_5 sp6_5 sp7_5 11.551961
Rsn6_5 sn6_5 sn7_5 11.551961
Rsp6_6 sp6_6 sp7_6 11.551961
Rsn6_6 sn6_6 sn7_6 11.551961
Rsp6_7 sp6_7 sp7_7 11.551961
Rsn6_7 sn6_7 sn7_7 11.551961
Rsp6_8 sp6_8 sp7_8 11.551961
Rsn6_8 sn6_8 sn7_8 11.551961
Rsp6_9 sp6_9 sp7_9 11.551961
Rsn6_9 sn6_9 sn7_9 11.551961
Rsp6_10 sp6_10 sp7_10 11.551961
Rsn6_10 sn6_10 sn7_10 11.551961
Rsp7_1 sp7_1 sp8_1 11.551961
Rsn7_1 sn7_1 sn8_1 11.551961
Rsp7_2 sp7_2 sp8_2 11.551961
Rsn7_2 sn7_2 sn8_2 11.551961
Rsp7_3 sp7_3 sp8_3 11.551961
Rsn7_3 sn7_3 sn8_3 11.551961
Rsp7_4 sp7_4 sp8_4 11.551961
Rsn7_4 sn7_4 sn8_4 11.551961
Rsp7_5 sp7_5 sp8_5 11.551961
Rsn7_5 sn7_5 sn8_5 11.551961
Rsp7_6 sp7_6 sp8_6 11.551961
Rsn7_6 sn7_6 sn8_6 11.551961
Rsp7_7 sp7_7 sp8_7 11.551961
Rsn7_7 sn7_7 sn8_7 11.551961
Rsp7_8 sp7_8 sp8_8 11.551961
Rsn7_8 sn7_8 sn8_8 11.551961
Rsp7_9 sp7_9 sp8_9 11.551961
Rsn7_9 sn7_9 sn8_9 11.551961
Rsp7_10 sp7_10 sp8_10 11.551961
Rsn7_10 sn7_10 sn8_10 11.551961
Rsp8_1 sp8_1 sp9_1 11.551961
Rsn8_1 sn8_1 sn9_1 11.551961
Rsp8_2 sp8_2 sp9_2 11.551961
Rsn8_2 sn8_2 sn9_2 11.551961
Rsp8_3 sp8_3 sp9_3 11.551961
Rsn8_3 sn8_3 sn9_3 11.551961
Rsp8_4 sp8_4 sp9_4 11.551961
Rsn8_4 sn8_4 sn9_4 11.551961
Rsp8_5 sp8_5 sp9_5 11.551961
Rsn8_5 sn8_5 sn9_5 11.551961
Rsp8_6 sp8_6 sp9_6 11.551961
Rsn8_6 sn8_6 sn9_6 11.551961
Rsp8_7 sp8_7 sp9_7 11.551961
Rsn8_7 sn8_7 sn9_7 11.551961
Rsp8_8 sp8_8 sp9_8 11.551961
Rsn8_8 sn8_8 sn9_8 11.551961
Rsp8_9 sp8_9 sp9_9 11.551961
Rsn8_9 sn8_9 sn9_9 11.551961
Rsp8_10 sp8_10 sp9_10 11.551961
Rsn8_10 sn8_10 sn9_10 11.551961
Rsp9_1 sp9_1 sp10_1 11.551961
Rsn9_1 sn9_1 sn10_1 11.551961
Rsp9_2 sp9_2 sp10_2 11.551961
Rsn9_2 sn9_2 sn10_2 11.551961
Rsp9_3 sp9_3 sp10_3 11.551961
Rsn9_3 sn9_3 sn10_3 11.551961
Rsp9_4 sp9_4 sp10_4 11.551961
Rsn9_4 sn9_4 sn10_4 11.551961
Rsp9_5 sp9_5 sp10_5 11.551961
Rsn9_5 sn9_5 sn10_5 11.551961
Rsp9_6 sp9_6 sp10_6 11.551961
Rsn9_6 sn9_6 sn10_6 11.551961
Rsp9_7 sp9_7 sp10_7 11.551961
Rsn9_7 sn9_7 sn10_7 11.551961
Rsp9_8 sp9_8 sp10_8 11.551961
Rsn9_8 sn9_8 sn10_8 11.551961
Rsp9_9 sp9_9 sp10_9 11.551961
Rsn9_9 sn9_9 sn10_9 11.551961
Rsp9_10 sp9_10 sp10_10 11.551961
Rsn9_10 sn9_10 sn10_10 11.551961
Rsp10_1 sp10_1 sp11_1 11.551961
Rsn10_1 sn10_1 sn11_1 11.551961
Rsp10_2 sp10_2 sp11_2 11.551961
Rsn10_2 sn10_2 sn11_2 11.551961
Rsp10_3 sp10_3 sp11_3 11.551961
Rsn10_3 sn10_3 sn11_3 11.551961
Rsp10_4 sp10_4 sp11_4 11.551961
Rsn10_4 sn10_4 sn11_4 11.551961
Rsp10_5 sp10_5 sp11_5 11.551961
Rsn10_5 sn10_5 sn11_5 11.551961
Rsp10_6 sp10_6 sp11_6 11.551961
Rsn10_6 sn10_6 sn11_6 11.551961
Rsp10_7 sp10_7 sp11_7 11.551961
Rsn10_7 sn10_7 sn11_7 11.551961
Rsp10_8 sp10_8 sp11_8 11.551961
Rsn10_8 sn10_8 sn11_8 11.551961
Rsp10_9 sp10_9 sp11_9 11.551961
Rsn10_9 sn10_9 sn11_9 11.551961
Rsp10_10 sp10_10 sp11_10 11.551961
Rsn10_10 sn10_10 sn11_10 11.551961
Rsp11_1 sp11_1 sp12_1 11.551961
Rsn11_1 sn11_1 sn12_1 11.551961
Rsp11_2 sp11_2 sp12_2 11.551961
Rsn11_2 sn11_2 sn12_2 11.551961
Rsp11_3 sp11_3 sp12_3 11.551961
Rsn11_3 sn11_3 sn12_3 11.551961
Rsp11_4 sp11_4 sp12_4 11.551961
Rsn11_4 sn11_4 sn12_4 11.551961
Rsp11_5 sp11_5 sp12_5 11.551961
Rsn11_5 sn11_5 sn12_5 11.551961
Rsp11_6 sp11_6 sp12_6 11.551961
Rsn11_6 sn11_6 sn12_6 11.551961
Rsp11_7 sp11_7 sp12_7 11.551961
Rsn11_7 sn11_7 sn12_7 11.551961
Rsp11_8 sp11_8 sp12_8 11.551961
Rsn11_8 sn11_8 sn12_8 11.551961
Rsp11_9 sp11_9 sp12_9 11.551961
Rsn11_9 sn11_9 sn12_9 11.551961
Rsp11_10 sp11_10 sp12_10 11.551961
Rsn11_10 sn11_10 sn12_10 11.551961
Rsp12_1 sp12_1 sp13_1 11.551961
Rsn12_1 sn12_1 sn13_1 11.551961
Rsp12_2 sp12_2 sp13_2 11.551961
Rsn12_2 sn12_2 sn13_2 11.551961
Rsp12_3 sp12_3 sp13_3 11.551961
Rsn12_3 sn12_3 sn13_3 11.551961
Rsp12_4 sp12_4 sp13_4 11.551961
Rsn12_4 sn12_4 sn13_4 11.551961
Rsp12_5 sp12_5 sp13_5 11.551961
Rsn12_5 sn12_5 sn13_5 11.551961
Rsp12_6 sp12_6 sp13_6 11.551961
Rsn12_6 sn12_6 sn13_6 11.551961
Rsp12_7 sp12_7 sp13_7 11.551961
Rsn12_7 sn12_7 sn13_7 11.551961
Rsp12_8 sp12_8 sp13_8 11.551961
Rsn12_8 sn12_8 sn13_8 11.551961
Rsp12_9 sp12_9 sp13_9 11.551961
Rsn12_9 sn12_9 sn13_9 11.551961
Rsp12_10 sp12_10 sp13_10 11.551961
Rsn12_10 sn12_10 sn13_10 11.551961
Rsp13_1 sp13_1 sp14_1 11.551961
Rsn13_1 sn13_1 sn14_1 11.551961
Rsp13_2 sp13_2 sp14_2 11.551961
Rsn13_2 sn13_2 sn14_2 11.551961
Rsp13_3 sp13_3 sp14_3 11.551961
Rsn13_3 sn13_3 sn14_3 11.551961
Rsp13_4 sp13_4 sp14_4 11.551961
Rsn13_4 sn13_4 sn14_4 11.551961
Rsp13_5 sp13_5 sp14_5 11.551961
Rsn13_5 sn13_5 sn14_5 11.551961
Rsp13_6 sp13_6 sp14_6 11.551961
Rsn13_6 sn13_6 sn14_6 11.551961
Rsp13_7 sp13_7 sp14_7 11.551961
Rsn13_7 sn13_7 sn14_7 11.551961
Rsp13_8 sp13_8 sp14_8 11.551961
Rsn13_8 sn13_8 sn14_8 11.551961
Rsp13_9 sp13_9 sp14_9 11.551961
Rsn13_9 sn13_9 sn14_9 11.551961
Rsp13_10 sp13_10 sp14_10 11.551961
Rsn13_10 sn13_10 sn14_10 11.551961
Rsp14_1 sp14_1 sp15_1 11.551961
Rsn14_1 sn14_1 sn15_1 11.551961
Rsp14_2 sp14_2 sp15_2 11.551961
Rsn14_2 sn14_2 sn15_2 11.551961
Rsp14_3 sp14_3 sp15_3 11.551961
Rsn14_3 sn14_3 sn15_3 11.551961
Rsp14_4 sp14_4 sp15_4 11.551961
Rsn14_4 sn14_4 sn15_4 11.551961
Rsp14_5 sp14_5 sp15_5 11.551961
Rsn14_5 sn14_5 sn15_5 11.551961
Rsp14_6 sp14_6 sp15_6 11.551961
Rsn14_6 sn14_6 sn15_6 11.551961
Rsp14_7 sp14_7 sp15_7 11.551961
Rsn14_7 sn14_7 sn15_7 11.551961
Rsp14_8 sp14_8 sp15_8 11.551961
Rsn14_8 sn14_8 sn15_8 11.551961
Rsp14_9 sp14_9 sp15_9 11.551961
Rsn14_9 sn14_9 sn15_9 11.551961
Rsp14_10 sp14_10 sp15_10 11.551961
Rsn14_10 sn14_10 sn15_10 11.551961
Rsp15_1 sp15_1 sp16_1 11.551961
Rsn15_1 sn15_1 sn16_1 11.551961
Rsp15_2 sp15_2 sp16_2 11.551961
Rsn15_2 sn15_2 sn16_2 11.551961
Rsp15_3 sp15_3 sp16_3 11.551961
Rsn15_3 sn15_3 sn16_3 11.551961
Rsp15_4 sp15_4 sp16_4 11.551961
Rsn15_4 sn15_4 sn16_4 11.551961
Rsp15_5 sp15_5 sp16_5 11.551961
Rsn15_5 sn15_5 sn16_5 11.551961
Rsp15_6 sp15_6 sp16_6 11.551961
Rsn15_6 sn15_6 sn16_6 11.551961
Rsp15_7 sp15_7 sp16_7 11.551961
Rsn15_7 sn15_7 sn16_7 11.551961
Rsp15_8 sp15_8 sp16_8 11.551961
Rsn15_8 sn15_8 sn16_8 11.551961
Rsp15_9 sp15_9 sp16_9 11.551961
Rsn15_9 sn15_9 sn16_9 11.551961
Rsp15_10 sp15_10 sp16_10 11.551961
Rsn15_10 sn15_10 sn16_10 11.551961
Rsp16_1 sp16_1 sp17_1 11.551961
Rsn16_1 sn16_1 sn17_1 11.551961
Rsp16_2 sp16_2 sp17_2 11.551961
Rsn16_2 sn16_2 sn17_2 11.551961
Rsp16_3 sp16_3 sp17_3 11.551961
Rsn16_3 sn16_3 sn17_3 11.551961
Rsp16_4 sp16_4 sp17_4 11.551961
Rsn16_4 sn16_4 sn17_4 11.551961
Rsp16_5 sp16_5 sp17_5 11.551961
Rsn16_5 sn16_5 sn17_5 11.551961
Rsp16_6 sp16_6 sp17_6 11.551961
Rsn16_6 sn16_6 sn17_6 11.551961
Rsp16_7 sp16_7 sp17_7 11.551961
Rsn16_7 sn16_7 sn17_7 11.551961
Rsp16_8 sp16_8 sp17_8 11.551961
Rsn16_8 sn16_8 sn17_8 11.551961
Rsp16_9 sp16_9 sp17_9 11.551961
Rsn16_9 sn16_9 sn17_9 11.551961
Rsp16_10 sp16_10 sp17_10 11.551961
Rsn16_10 sn16_10 sn17_10 11.551961
Rsp17_1 sp17_1 sp18_1 11.551961
Rsn17_1 sn17_1 sn18_1 11.551961
Rsp17_2 sp17_2 sp18_2 11.551961
Rsn17_2 sn17_2 sn18_2 11.551961
Rsp17_3 sp17_3 sp18_3 11.551961
Rsn17_3 sn17_3 sn18_3 11.551961
Rsp17_4 sp17_4 sp18_4 11.551961
Rsn17_4 sn17_4 sn18_4 11.551961
Rsp17_5 sp17_5 sp18_5 11.551961
Rsn17_5 sn17_5 sn18_5 11.551961
Rsp17_6 sp17_6 sp18_6 11.551961
Rsn17_6 sn17_6 sn18_6 11.551961
Rsp17_7 sp17_7 sp18_7 11.551961
Rsn17_7 sn17_7 sn18_7 11.551961
Rsp17_8 sp17_8 sp18_8 11.551961
Rsn17_8 sn17_8 sn18_8 11.551961
Rsp17_9 sp17_9 sp18_9 11.551961
Rsn17_9 sn17_9 sn18_9 11.551961
Rsp17_10 sp17_10 sp18_10 11.551961
Rsn17_10 sn17_10 sn18_10 11.551961
Rsp18_1 sp18_1 sp19_1 11.551961
Rsn18_1 sn18_1 sn19_1 11.551961
Rsp18_2 sp18_2 sp19_2 11.551961
Rsn18_2 sn18_2 sn19_2 11.551961
Rsp18_3 sp18_3 sp19_3 11.551961
Rsn18_3 sn18_3 sn19_3 11.551961
Rsp18_4 sp18_4 sp19_4 11.551961
Rsn18_4 sn18_4 sn19_4 11.551961
Rsp18_5 sp18_5 sp19_5 11.551961
Rsn18_5 sn18_5 sn19_5 11.551961
Rsp18_6 sp18_6 sp19_6 11.551961
Rsn18_6 sn18_6 sn19_6 11.551961
Rsp18_7 sp18_7 sp19_7 11.551961
Rsn18_7 sn18_7 sn19_7 11.551961
Rsp18_8 sp18_8 sp19_8 11.551961
Rsn18_8 sn18_8 sn19_8 11.551961
Rsp18_9 sp18_9 sp19_9 11.551961
Rsn18_9 sn18_9 sn19_9 11.551961
Rsp18_10 sp18_10 sp19_10 11.551961
Rsn18_10 sn18_10 sn19_10 11.551961
Rsp19_1 sp19_1 sp20_1 11.551961
Rsn19_1 sn19_1 sn20_1 11.551961
Rsp19_2 sp19_2 sp20_2 11.551961
Rsn19_2 sn19_2 sn20_2 11.551961
Rsp19_3 sp19_3 sp20_3 11.551961
Rsn19_3 sn19_3 sn20_3 11.551961
Rsp19_4 sp19_4 sp20_4 11.551961
Rsn19_4 sn19_4 sn20_4 11.551961
Rsp19_5 sp19_5 sp20_5 11.551961
Rsn19_5 sn19_5 sn20_5 11.551961
Rsp19_6 sp19_6 sp20_6 11.551961
Rsn19_6 sn19_6 sn20_6 11.551961
Rsp19_7 sp19_7 sp20_7 11.551961
Rsn19_7 sn19_7 sn20_7 11.551961
Rsp19_8 sp19_8 sp20_8 11.551961
Rsn19_8 sn19_8 sn20_8 11.551961
Rsp19_9 sp19_9 sp20_9 11.551961
Rsn19_9 sn19_9 sn20_9 11.551961
Rsp19_10 sp19_10 sp20_10 11.551961
Rsn19_10 sn19_10 sn20_10 11.551961
Rsp20_1 sp20_1 sp21_1 11.551961
Rsn20_1 sn20_1 sn21_1 11.551961
Rsp20_2 sp20_2 sp21_2 11.551961
Rsn20_2 sn20_2 sn21_2 11.551961
Rsp20_3 sp20_3 sp21_3 11.551961
Rsn20_3 sn20_3 sn21_3 11.551961
Rsp20_4 sp20_4 sp21_4 11.551961
Rsn20_4 sn20_4 sn21_4 11.551961
Rsp20_5 sp20_5 sp21_5 11.551961
Rsn20_5 sn20_5 sn21_5 11.551961
Rsp20_6 sp20_6 sp21_6 11.551961
Rsn20_6 sn20_6 sn21_6 11.551961
Rsp20_7 sp20_7 sp21_7 11.551961
Rsn20_7 sn20_7 sn21_7 11.551961
Rsp20_8 sp20_8 sp21_8 11.551961
Rsn20_8 sn20_8 sn21_8 11.551961
Rsp20_9 sp20_9 sp21_9 11.551961
Rsn20_9 sn20_9 sn21_9 11.551961
Rsp20_10 sp20_10 sp21_10 11.551961
Rsn20_10 sn20_10 sn21_10 11.551961
Rsp21_1 sp21_1 sp22_1 11.551961
Rsn21_1 sn21_1 sn22_1 11.551961
Rsp21_2 sp21_2 sp22_2 11.551961
Rsn21_2 sn21_2 sn22_2 11.551961
Rsp21_3 sp21_3 sp22_3 11.551961
Rsn21_3 sn21_3 sn22_3 11.551961
Rsp21_4 sp21_4 sp22_4 11.551961
Rsn21_4 sn21_4 sn22_4 11.551961
Rsp21_5 sp21_5 sp22_5 11.551961
Rsn21_5 sn21_5 sn22_5 11.551961
Rsp21_6 sp21_6 sp22_6 11.551961
Rsn21_6 sn21_6 sn22_6 11.551961
Rsp21_7 sp21_7 sp22_7 11.551961
Rsn21_7 sn21_7 sn22_7 11.551961
Rsp21_8 sp21_8 sp22_8 11.551961
Rsn21_8 sn21_8 sn22_8 11.551961
Rsp21_9 sp21_9 sp22_9 11.551961
Rsn21_9 sn21_9 sn22_9 11.551961
Rsp21_10 sp21_10 sp22_10 11.551961
Rsn21_10 sn21_10 sn22_10 11.551961
Rsp22_1 sp22_1 sp23_1 11.551961
Rsn22_1 sn22_1 sn23_1 11.551961
Rsp22_2 sp22_2 sp23_2 11.551961
Rsn22_2 sn22_2 sn23_2 11.551961
Rsp22_3 sp22_3 sp23_3 11.551961
Rsn22_3 sn22_3 sn23_3 11.551961
Rsp22_4 sp22_4 sp23_4 11.551961
Rsn22_4 sn22_4 sn23_4 11.551961
Rsp22_5 sp22_5 sp23_5 11.551961
Rsn22_5 sn22_5 sn23_5 11.551961
Rsp22_6 sp22_6 sp23_6 11.551961
Rsn22_6 sn22_6 sn23_6 11.551961
Rsp22_7 sp22_7 sp23_7 11.551961
Rsn22_7 sn22_7 sn23_7 11.551961
Rsp22_8 sp22_8 sp23_8 11.551961
Rsn22_8 sn22_8 sn23_8 11.551961
Rsp22_9 sp22_9 sp23_9 11.551961
Rsn22_9 sn22_9 sn23_9 11.551961
Rsp22_10 sp22_10 sp23_10 11.551961
Rsn22_10 sn22_10 sn23_10 11.551961
Rsp23_1 sp23_1 sp24_1 11.551961
Rsn23_1 sn23_1 sn24_1 11.551961
Rsp23_2 sp23_2 sp24_2 11.551961
Rsn23_2 sn23_2 sn24_2 11.551961
Rsp23_3 sp23_3 sp24_3 11.551961
Rsn23_3 sn23_3 sn24_3 11.551961
Rsp23_4 sp23_4 sp24_4 11.551961
Rsn23_4 sn23_4 sn24_4 11.551961
Rsp23_5 sp23_5 sp24_5 11.551961
Rsn23_5 sn23_5 sn24_5 11.551961
Rsp23_6 sp23_6 sp24_6 11.551961
Rsn23_6 sn23_6 sn24_6 11.551961
Rsp23_7 sp23_7 sp24_7 11.551961
Rsn23_7 sn23_7 sn24_7 11.551961
Rsp23_8 sp23_8 sp24_8 11.551961
Rsn23_8 sn23_8 sn24_8 11.551961
Rsp23_9 sp23_9 sp24_9 11.551961
Rsn23_9 sn23_9 sn24_9 11.551961
Rsp23_10 sp23_10 sp24_10 11.551961
Rsn23_10 sn23_10 sn24_10 11.551961
Rsp24_1 sp24_1 sp25_1 11.551961
Rsn24_1 sn24_1 sn25_1 11.551961
Rsp24_2 sp24_2 sp25_2 11.551961
Rsn24_2 sn24_2 sn25_2 11.551961
Rsp24_3 sp24_3 sp25_3 11.551961
Rsn24_3 sn24_3 sn25_3 11.551961
Rsp24_4 sp24_4 sp25_4 11.551961
Rsn24_4 sn24_4 sn25_4 11.551961
Rsp24_5 sp24_5 sp25_5 11.551961
Rsn24_5 sn24_5 sn25_5 11.551961
Rsp24_6 sp24_6 sp25_6 11.551961
Rsn24_6 sn24_6 sn25_6 11.551961
Rsp24_7 sp24_7 sp25_7 11.551961
Rsn24_7 sn24_7 sn25_7 11.551961
Rsp24_8 sp24_8 sp25_8 11.551961
Rsn24_8 sn24_8 sn25_8 11.551961
Rsp24_9 sp24_9 sp25_9 11.551961
Rsn24_9 sn24_9 sn25_9 11.551961
Rsp24_10 sp24_10 sp25_10 11.551961
Rsn24_10 sn24_10 sn25_10 11.551961
Rsp25_1 sp25_1 sp26_1 11.551961
Rsn25_1 sn25_1 sn26_1 11.551961
Rsp25_2 sp25_2 sp26_2 11.551961
Rsn25_2 sn25_2 sn26_2 11.551961
Rsp25_3 sp25_3 sp26_3 11.551961
Rsn25_3 sn25_3 sn26_3 11.551961
Rsp25_4 sp25_4 sp26_4 11.551961
Rsn25_4 sn25_4 sn26_4 11.551961
Rsp25_5 sp25_5 sp26_5 11.551961
Rsn25_5 sn25_5 sn26_5 11.551961
Rsp25_6 sp25_6 sp26_6 11.551961
Rsn25_6 sn25_6 sn26_6 11.551961
Rsp25_7 sp25_7 sp26_7 11.551961
Rsn25_7 sn25_7 sn26_7 11.551961
Rsp25_8 sp25_8 sp26_8 11.551961
Rsn25_8 sn25_8 sn26_8 11.551961
Rsp25_9 sp25_9 sp26_9 11.551961
Rsn25_9 sn25_9 sn26_9 11.551961
Rsp25_10 sp25_10 sp26_10 11.551961
Rsn25_10 sn25_10 sn26_10 11.551961
Rsp26_1 sp26_1 sp27_1 11.551961
Rsn26_1 sn26_1 sn27_1 11.551961
Rsp26_2 sp26_2 sp27_2 11.551961
Rsn26_2 sn26_2 sn27_2 11.551961
Rsp26_3 sp26_3 sp27_3 11.551961
Rsn26_3 sn26_3 sn27_3 11.551961
Rsp26_4 sp26_4 sp27_4 11.551961
Rsn26_4 sn26_4 sn27_4 11.551961
Rsp26_5 sp26_5 sp27_5 11.551961
Rsn26_5 sn26_5 sn27_5 11.551961
Rsp26_6 sp26_6 sp27_6 11.551961
Rsn26_6 sn26_6 sn27_6 11.551961
Rsp26_7 sp26_7 sp27_7 11.551961
Rsn26_7 sn26_7 sn27_7 11.551961
Rsp26_8 sp26_8 sp27_8 11.551961
Rsn26_8 sn26_8 sn27_8 11.551961
Rsp26_9 sp26_9 sp27_9 11.551961
Rsn26_9 sn26_9 sn27_9 11.551961
Rsp26_10 sp26_10 sp27_10 11.551961
Rsn26_10 sn26_10 sn27_10 11.551961
Rsp27_1 sp27_1 sp28_1 11.551961
Rsn27_1 sn27_1 sn28_1 11.551961
Rsp27_2 sp27_2 sp28_2 11.551961
Rsn27_2 sn27_2 sn28_2 11.551961
Rsp27_3 sp27_3 sp28_3 11.551961
Rsn27_3 sn27_3 sn28_3 11.551961
Rsp27_4 sp27_4 sp28_4 11.551961
Rsn27_4 sn27_4 sn28_4 11.551961
Rsp27_5 sp27_5 sp28_5 11.551961
Rsn27_5 sn27_5 sn28_5 11.551961
Rsp27_6 sp27_6 sp28_6 11.551961
Rsn27_6 sn27_6 sn28_6 11.551961
Rsp27_7 sp27_7 sp28_7 11.551961
Rsn27_7 sn27_7 sn28_7 11.551961
Rsp27_8 sp27_8 sp28_8 11.551961
Rsn27_8 sn27_8 sn28_8 11.551961
Rsp27_9 sp27_9 sp28_9 11.551961
Rsn27_9 sn27_9 sn28_9 11.551961
Rsp27_10 sp27_10 sp28_10 11.551961
Rsn27_10 sn27_10 sn28_10 11.551961
Rsp28_1 sp28_1 sp29_1 11.551961
Rsn28_1 sn28_1 sn29_1 11.551961
Rsp28_2 sp28_2 sp29_2 11.551961
Rsn28_2 sn28_2 sn29_2 11.551961
Rsp28_3 sp28_3 sp29_3 11.551961
Rsn28_3 sn28_3 sn29_3 11.551961
Rsp28_4 sp28_4 sp29_4 11.551961
Rsn28_4 sn28_4 sn29_4 11.551961
Rsp28_5 sp28_5 sp29_5 11.551961
Rsn28_5 sn28_5 sn29_5 11.551961
Rsp28_6 sp28_6 sp29_6 11.551961
Rsn28_6 sn28_6 sn29_6 11.551961
Rsp28_7 sp28_7 sp29_7 11.551961
Rsn28_7 sn28_7 sn29_7 11.551961
Rsp28_8 sp28_8 sp29_8 11.551961
Rsn28_8 sn28_8 sn29_8 11.551961
Rsp28_9 sp28_9 sp29_9 11.551961
Rsn28_9 sn28_9 sn29_9 11.551961
Rsp28_10 sp28_10 sp29_10 11.551961
Rsn28_10 sn28_10 sn29_10 11.551961
Rsp29_1 sp29_1 sp1_p1 11.551961
Rsn29_1 sn29_1 sn1_p1 11.551961
Rsp29_2 sp29_2 sp2_p1 11.551961
Rsn29_2 sn29_2 sn2_p1 11.551961
Rsp29_3 sp29_3 sp3_p1 11.551961
Rsn29_3 sn29_3 sn3_p1 11.551961
Rsp29_4 sp29_4 sp4_p1 11.551961
Rsn29_4 sn29_4 sn4_p1 11.551961
Rsp29_5 sp29_5 sp5_p1 11.551961
Rsn29_5 sn29_5 sn5_p1 11.551961
Rsp29_6 sp29_6 sp6_p1 11.551961
Rsn29_6 sn29_6 sn6_p1 11.551961
Rsp29_7 sp29_7 sp7_p1 11.551961
Rsn29_7 sn29_7 sn7_p1 11.551961
Rsp29_8 sp29_8 sp8_p1 11.551961
Rsn29_8 sn29_8 sn8_p1 11.551961
Rsp29_9 sp29_9 sp9_p1 11.551961
Rsn29_9 sn29_9 sn9_p1 11.551961
Rsp29_10 sp29_10 sp10_p1 11.551961
Rsn29_10 sn29_10 sn10_p1 11.551961
Rsp30_1 sp30_1 sp31_1 11.551961
Rsn30_1 sn30_1 sn31_1 11.551961
Rsp30_2 sp30_2 sp31_2 11.551961
Rsn30_2 sn30_2 sn31_2 11.551961
Rsp30_3 sp30_3 sp31_3 11.551961
Rsn30_3 sn30_3 sn31_3 11.551961
Rsp30_4 sp30_4 sp31_4 11.551961
Rsn30_4 sn30_4 sn31_4 11.551961
Rsp30_5 sp30_5 sp31_5 11.551961
Rsn30_5 sn30_5 sn31_5 11.551961
Rsp30_6 sp30_6 sp31_6 11.551961
Rsn30_6 sn30_6 sn31_6 11.551961
Rsp30_7 sp30_7 sp31_7 11.551961
Rsn30_7 sn30_7 sn31_7 11.551961
Rsp30_8 sp30_8 sp31_8 11.551961
Rsn30_8 sn30_8 sn31_8 11.551961
Rsp30_9 sp30_9 sp31_9 11.551961
Rsn30_9 sn30_9 sn31_9 11.551961
Rsp30_10 sp30_10 sp31_10 11.551961
Rsn30_10 sn30_10 sn31_10 11.551961
Rsp31_1 sp31_1 sp32_1 11.551961
Rsn31_1 sn31_1 sn32_1 11.551961
Rsp31_2 sp31_2 sp32_2 11.551961
Rsn31_2 sn31_2 sn32_2 11.551961
Rsp31_3 sp31_3 sp32_3 11.551961
Rsn31_3 sn31_3 sn32_3 11.551961
Rsp31_4 sp31_4 sp32_4 11.551961
Rsn31_4 sn31_4 sn32_4 11.551961
Rsp31_5 sp31_5 sp32_5 11.551961
Rsn31_5 sn31_5 sn32_5 11.551961
Rsp31_6 sp31_6 sp32_6 11.551961
Rsn31_6 sn31_6 sn32_6 11.551961
Rsp31_7 sp31_7 sp32_7 11.551961
Rsn31_7 sn31_7 sn32_7 11.551961
Rsp31_8 sp31_8 sp32_8 11.551961
Rsn31_8 sn31_8 sn32_8 11.551961
Rsp31_9 sp31_9 sp32_9 11.551961
Rsn31_9 sn31_9 sn32_9 11.551961
Rsp31_10 sp31_10 sp32_10 11.551961
Rsn31_10 sn31_10 sn32_10 11.551961
Rsp32_1 sp32_1 sp33_1 11.551961
Rsn32_1 sn32_1 sn33_1 11.551961
Rsp32_2 sp32_2 sp33_2 11.551961
Rsn32_2 sn32_2 sn33_2 11.551961
Rsp32_3 sp32_3 sp33_3 11.551961
Rsn32_3 sn32_3 sn33_3 11.551961
Rsp32_4 sp32_4 sp33_4 11.551961
Rsn32_4 sn32_4 sn33_4 11.551961
Rsp32_5 sp32_5 sp33_5 11.551961
Rsn32_5 sn32_5 sn33_5 11.551961
Rsp32_6 sp32_6 sp33_6 11.551961
Rsn32_6 sn32_6 sn33_6 11.551961
Rsp32_7 sp32_7 sp33_7 11.551961
Rsn32_7 sn32_7 sn33_7 11.551961
Rsp32_8 sp32_8 sp33_8 11.551961
Rsn32_8 sn32_8 sn33_8 11.551961
Rsp32_9 sp32_9 sp33_9 11.551961
Rsn32_9 sn32_9 sn33_9 11.551961
Rsp32_10 sp32_10 sp33_10 11.551961
Rsn32_10 sn32_10 sn33_10 11.551961
Rsp33_1 sp33_1 sp34_1 11.551961
Rsn33_1 sn33_1 sn34_1 11.551961
Rsp33_2 sp33_2 sp34_2 11.551961
Rsn33_2 sn33_2 sn34_2 11.551961
Rsp33_3 sp33_3 sp34_3 11.551961
Rsn33_3 sn33_3 sn34_3 11.551961
Rsp33_4 sp33_4 sp34_4 11.551961
Rsn33_4 sn33_4 sn34_4 11.551961
Rsp33_5 sp33_5 sp34_5 11.551961
Rsn33_5 sn33_5 sn34_5 11.551961
Rsp33_6 sp33_6 sp34_6 11.551961
Rsn33_6 sn33_6 sn34_6 11.551961
Rsp33_7 sp33_7 sp34_7 11.551961
Rsn33_7 sn33_7 sn34_7 11.551961
Rsp33_8 sp33_8 sp34_8 11.551961
Rsn33_8 sn33_8 sn34_8 11.551961
Rsp33_9 sp33_9 sp34_9 11.551961
Rsn33_9 sn33_9 sn34_9 11.551961
Rsp33_10 sp33_10 sp34_10 11.551961
Rsn33_10 sn33_10 sn34_10 11.551961
Rsp34_1 sp34_1 sp35_1 11.551961
Rsn34_1 sn34_1 sn35_1 11.551961
Rsp34_2 sp34_2 sp35_2 11.551961
Rsn34_2 sn34_2 sn35_2 11.551961
Rsp34_3 sp34_3 sp35_3 11.551961
Rsn34_3 sn34_3 sn35_3 11.551961
Rsp34_4 sp34_4 sp35_4 11.551961
Rsn34_4 sn34_4 sn35_4 11.551961
Rsp34_5 sp34_5 sp35_5 11.551961
Rsn34_5 sn34_5 sn35_5 11.551961
Rsp34_6 sp34_6 sp35_6 11.551961
Rsn34_6 sn34_6 sn35_6 11.551961
Rsp34_7 sp34_7 sp35_7 11.551961
Rsn34_7 sn34_7 sn35_7 11.551961
Rsp34_8 sp34_8 sp35_8 11.551961
Rsn34_8 sn34_8 sn35_8 11.551961
Rsp34_9 sp34_9 sp35_9 11.551961
Rsn34_9 sn34_9 sn35_9 11.551961
Rsp34_10 sp34_10 sp35_10 11.551961
Rsn34_10 sn34_10 sn35_10 11.551961
Rsp35_1 sp35_1 sp36_1 11.551961
Rsn35_1 sn35_1 sn36_1 11.551961
Rsp35_2 sp35_2 sp36_2 11.551961
Rsn35_2 sn35_2 sn36_2 11.551961
Rsp35_3 sp35_3 sp36_3 11.551961
Rsn35_3 sn35_3 sn36_3 11.551961
Rsp35_4 sp35_4 sp36_4 11.551961
Rsn35_4 sn35_4 sn36_4 11.551961
Rsp35_5 sp35_5 sp36_5 11.551961
Rsn35_5 sn35_5 sn36_5 11.551961
Rsp35_6 sp35_6 sp36_6 11.551961
Rsn35_6 sn35_6 sn36_6 11.551961
Rsp35_7 sp35_7 sp36_7 11.551961
Rsn35_7 sn35_7 sn36_7 11.551961
Rsp35_8 sp35_8 sp36_8 11.551961
Rsn35_8 sn35_8 sn36_8 11.551961
Rsp35_9 sp35_9 sp36_9 11.551961
Rsn35_9 sn35_9 sn36_9 11.551961
Rsp35_10 sp35_10 sp36_10 11.551961
Rsn35_10 sn35_10 sn36_10 11.551961
Rsp36_1 sp36_1 sp37_1 11.551961
Rsn36_1 sn36_1 sn37_1 11.551961
Rsp36_2 sp36_2 sp37_2 11.551961
Rsn36_2 sn36_2 sn37_2 11.551961
Rsp36_3 sp36_3 sp37_3 11.551961
Rsn36_3 sn36_3 sn37_3 11.551961
Rsp36_4 sp36_4 sp37_4 11.551961
Rsn36_4 sn36_4 sn37_4 11.551961
Rsp36_5 sp36_5 sp37_5 11.551961
Rsn36_5 sn36_5 sn37_5 11.551961
Rsp36_6 sp36_6 sp37_6 11.551961
Rsn36_6 sn36_6 sn37_6 11.551961
Rsp36_7 sp36_7 sp37_7 11.551961
Rsn36_7 sn36_7 sn37_7 11.551961
Rsp36_8 sp36_8 sp37_8 11.551961
Rsn36_8 sn36_8 sn37_8 11.551961
Rsp36_9 sp36_9 sp37_9 11.551961
Rsn36_9 sn36_9 sn37_9 11.551961
Rsp36_10 sp36_10 sp37_10 11.551961
Rsn36_10 sn36_10 sn37_10 11.551961
Rsp37_1 sp37_1 sp38_1 11.551961
Rsn37_1 sn37_1 sn38_1 11.551961
Rsp37_2 sp37_2 sp38_2 11.551961
Rsn37_2 sn37_2 sn38_2 11.551961
Rsp37_3 sp37_3 sp38_3 11.551961
Rsn37_3 sn37_3 sn38_3 11.551961
Rsp37_4 sp37_4 sp38_4 11.551961
Rsn37_4 sn37_4 sn38_4 11.551961
Rsp37_5 sp37_5 sp38_5 11.551961
Rsn37_5 sn37_5 sn38_5 11.551961
Rsp37_6 sp37_6 sp38_6 11.551961
Rsn37_6 sn37_6 sn38_6 11.551961
Rsp37_7 sp37_7 sp38_7 11.551961
Rsn37_7 sn37_7 sn38_7 11.551961
Rsp37_8 sp37_8 sp38_8 11.551961
Rsn37_8 sn37_8 sn38_8 11.551961
Rsp37_9 sp37_9 sp38_9 11.551961
Rsn37_9 sn37_9 sn38_9 11.551961
Rsp37_10 sp37_10 sp38_10 11.551961
Rsn37_10 sn37_10 sn38_10 11.551961
Rsp38_1 sp38_1 sp39_1 11.551961
Rsn38_1 sn38_1 sn39_1 11.551961
Rsp38_2 sp38_2 sp39_2 11.551961
Rsn38_2 sn38_2 sn39_2 11.551961
Rsp38_3 sp38_3 sp39_3 11.551961
Rsn38_3 sn38_3 sn39_3 11.551961
Rsp38_4 sp38_4 sp39_4 11.551961
Rsn38_4 sn38_4 sn39_4 11.551961
Rsp38_5 sp38_5 sp39_5 11.551961
Rsn38_5 sn38_5 sn39_5 11.551961
Rsp38_6 sp38_6 sp39_6 11.551961
Rsn38_6 sn38_6 sn39_6 11.551961
Rsp38_7 sp38_7 sp39_7 11.551961
Rsn38_7 sn38_7 sn39_7 11.551961
Rsp38_8 sp38_8 sp39_8 11.551961
Rsn38_8 sn38_8 sn39_8 11.551961
Rsp38_9 sp38_9 sp39_9 11.551961
Rsn38_9 sn38_9 sn39_9 11.551961
Rsp38_10 sp38_10 sp39_10 11.551961
Rsn38_10 sn38_10 sn39_10 11.551961
Rsp39_1 sp39_1 sp40_1 11.551961
Rsn39_1 sn39_1 sn40_1 11.551961
Rsp39_2 sp39_2 sp40_2 11.551961
Rsn39_2 sn39_2 sn40_2 11.551961
Rsp39_3 sp39_3 sp40_3 11.551961
Rsn39_3 sn39_3 sn40_3 11.551961
Rsp39_4 sp39_4 sp40_4 11.551961
Rsn39_4 sn39_4 sn40_4 11.551961
Rsp39_5 sp39_5 sp40_5 11.551961
Rsn39_5 sn39_5 sn40_5 11.551961
Rsp39_6 sp39_6 sp40_6 11.551961
Rsn39_6 sn39_6 sn40_6 11.551961
Rsp39_7 sp39_7 sp40_7 11.551961
Rsn39_7 sn39_7 sn40_7 11.551961
Rsp39_8 sp39_8 sp40_8 11.551961
Rsn39_8 sn39_8 sn40_8 11.551961
Rsp39_9 sp39_9 sp40_9 11.551961
Rsn39_9 sn39_9 sn40_9 11.551961
Rsp39_10 sp39_10 sp40_10 11.551961
Rsn39_10 sn39_10 sn40_10 11.551961
Rsp40_1 sp40_1 sp41_1 11.551961
Rsn40_1 sn40_1 sn41_1 11.551961
Rsp40_2 sp40_2 sp41_2 11.551961
Rsn40_2 sn40_2 sn41_2 11.551961
Rsp40_3 sp40_3 sp41_3 11.551961
Rsn40_3 sn40_3 sn41_3 11.551961
Rsp40_4 sp40_4 sp41_4 11.551961
Rsn40_4 sn40_4 sn41_4 11.551961
Rsp40_5 sp40_5 sp41_5 11.551961
Rsn40_5 sn40_5 sn41_5 11.551961
Rsp40_6 sp40_6 sp41_6 11.551961
Rsn40_6 sn40_6 sn41_6 11.551961
Rsp40_7 sp40_7 sp41_7 11.551961
Rsn40_7 sn40_7 sn41_7 11.551961
Rsp40_8 sp40_8 sp41_8 11.551961
Rsn40_8 sn40_8 sn41_8 11.551961
Rsp40_9 sp40_9 sp41_9 11.551961
Rsn40_9 sn40_9 sn41_9 11.551961
Rsp40_10 sp40_10 sp41_10 11.551961
Rsn40_10 sn40_10 sn41_10 11.551961
Rsp41_1 sp41_1 sp42_1 11.551961
Rsn41_1 sn41_1 sn42_1 11.551961
Rsp41_2 sp41_2 sp42_2 11.551961
Rsn41_2 sn41_2 sn42_2 11.551961
Rsp41_3 sp41_3 sp42_3 11.551961
Rsn41_3 sn41_3 sn42_3 11.551961
Rsp41_4 sp41_4 sp42_4 11.551961
Rsn41_4 sn41_4 sn42_4 11.551961
Rsp41_5 sp41_5 sp42_5 11.551961
Rsn41_5 sn41_5 sn42_5 11.551961
Rsp41_6 sp41_6 sp42_6 11.551961
Rsn41_6 sn41_6 sn42_6 11.551961
Rsp41_7 sp41_7 sp42_7 11.551961
Rsn41_7 sn41_7 sn42_7 11.551961
Rsp41_8 sp41_8 sp42_8 11.551961
Rsn41_8 sn41_8 sn42_8 11.551961
Rsp41_9 sp41_9 sp42_9 11.551961
Rsn41_9 sn41_9 sn42_9 11.551961
Rsp41_10 sp41_10 sp42_10 11.551961
Rsn41_10 sn41_10 sn42_10 11.551961
Rsp42_1 sp42_1 sp43_1 11.551961
Rsn42_1 sn42_1 sn43_1 11.551961
Rsp42_2 sp42_2 sp43_2 11.551961
Rsn42_2 sn42_2 sn43_2 11.551961
Rsp42_3 sp42_3 sp43_3 11.551961
Rsn42_3 sn42_3 sn43_3 11.551961
Rsp42_4 sp42_4 sp43_4 11.551961
Rsn42_4 sn42_4 sn43_4 11.551961
Rsp42_5 sp42_5 sp43_5 11.551961
Rsn42_5 sn42_5 sn43_5 11.551961
Rsp42_6 sp42_6 sp43_6 11.551961
Rsn42_6 sn42_6 sn43_6 11.551961
Rsp42_7 sp42_7 sp43_7 11.551961
Rsn42_7 sn42_7 sn43_7 11.551961
Rsp42_8 sp42_8 sp43_8 11.551961
Rsn42_8 sn42_8 sn43_8 11.551961
Rsp42_9 sp42_9 sp43_9 11.551961
Rsn42_9 sn42_9 sn43_9 11.551961
Rsp42_10 sp42_10 sp43_10 11.551961
Rsn42_10 sn42_10 sn43_10 11.551961
Rsp43_1 sp43_1 sp44_1 11.551961
Rsn43_1 sn43_1 sn44_1 11.551961
Rsp43_2 sp43_2 sp44_2 11.551961
Rsn43_2 sn43_2 sn44_2 11.551961
Rsp43_3 sp43_3 sp44_3 11.551961
Rsn43_3 sn43_3 sn44_3 11.551961
Rsp43_4 sp43_4 sp44_4 11.551961
Rsn43_4 sn43_4 sn44_4 11.551961
Rsp43_5 sp43_5 sp44_5 11.551961
Rsn43_5 sn43_5 sn44_5 11.551961
Rsp43_6 sp43_6 sp44_6 11.551961
Rsn43_6 sn43_6 sn44_6 11.551961
Rsp43_7 sp43_7 sp44_7 11.551961
Rsn43_7 sn43_7 sn44_7 11.551961
Rsp43_8 sp43_8 sp44_8 11.551961
Rsn43_8 sn43_8 sn44_8 11.551961
Rsp43_9 sp43_9 sp44_9 11.551961
Rsn43_9 sn43_9 sn44_9 11.551961
Rsp43_10 sp43_10 sp44_10 11.551961
Rsn43_10 sn43_10 sn44_10 11.551961
Rsp44_1 sp44_1 sp45_1 11.551961
Rsn44_1 sn44_1 sn45_1 11.551961
Rsp44_2 sp44_2 sp45_2 11.551961
Rsn44_2 sn44_2 sn45_2 11.551961
Rsp44_3 sp44_3 sp45_3 11.551961
Rsn44_3 sn44_3 sn45_3 11.551961
Rsp44_4 sp44_4 sp45_4 11.551961
Rsn44_4 sn44_4 sn45_4 11.551961
Rsp44_5 sp44_5 sp45_5 11.551961
Rsn44_5 sn44_5 sn45_5 11.551961
Rsp44_6 sp44_6 sp45_6 11.551961
Rsn44_6 sn44_6 sn45_6 11.551961
Rsp44_7 sp44_7 sp45_7 11.551961
Rsn44_7 sn44_7 sn45_7 11.551961
Rsp44_8 sp44_8 sp45_8 11.551961
Rsn44_8 sn44_8 sn45_8 11.551961
Rsp44_9 sp44_9 sp45_9 11.551961
Rsn44_9 sn44_9 sn45_9 11.551961
Rsp44_10 sp44_10 sp45_10 11.551961
Rsn44_10 sn44_10 sn45_10 11.551961
Rsp45_1 sp45_1 sp46_1 11.551961
Rsn45_1 sn45_1 sn46_1 11.551961
Rsp45_2 sp45_2 sp46_2 11.551961
Rsn45_2 sn45_2 sn46_2 11.551961
Rsp45_3 sp45_3 sp46_3 11.551961
Rsn45_3 sn45_3 sn46_3 11.551961
Rsp45_4 sp45_4 sp46_4 11.551961
Rsn45_4 sn45_4 sn46_4 11.551961
Rsp45_5 sp45_5 sp46_5 11.551961
Rsn45_5 sn45_5 sn46_5 11.551961
Rsp45_6 sp45_6 sp46_6 11.551961
Rsn45_6 sn45_6 sn46_6 11.551961
Rsp45_7 sp45_7 sp46_7 11.551961
Rsn45_7 sn45_7 sn46_7 11.551961
Rsp45_8 sp45_8 sp46_8 11.551961
Rsn45_8 sn45_8 sn46_8 11.551961
Rsp45_9 sp45_9 sp46_9 11.551961
Rsn45_9 sn45_9 sn46_9 11.551961
Rsp45_10 sp45_10 sp46_10 11.551961
Rsn45_10 sn45_10 sn46_10 11.551961
Rsp46_1 sp46_1 sp47_1 11.551961
Rsn46_1 sn46_1 sn47_1 11.551961
Rsp46_2 sp46_2 sp47_2 11.551961
Rsn46_2 sn46_2 sn47_2 11.551961
Rsp46_3 sp46_3 sp47_3 11.551961
Rsn46_3 sn46_3 sn47_3 11.551961
Rsp46_4 sp46_4 sp47_4 11.551961
Rsn46_4 sn46_4 sn47_4 11.551961
Rsp46_5 sp46_5 sp47_5 11.551961
Rsn46_5 sn46_5 sn47_5 11.551961
Rsp46_6 sp46_6 sp47_6 11.551961
Rsn46_6 sn46_6 sn47_6 11.551961
Rsp46_7 sp46_7 sp47_7 11.551961
Rsn46_7 sn46_7 sn47_7 11.551961
Rsp46_8 sp46_8 sp47_8 11.551961
Rsn46_8 sn46_8 sn47_8 11.551961
Rsp46_9 sp46_9 sp47_9 11.551961
Rsn46_9 sn46_9 sn47_9 11.551961
Rsp46_10 sp46_10 sp47_10 11.551961
Rsn46_10 sn46_10 sn47_10 11.551961
Rsp47_1 sp47_1 sp48_1 11.551961
Rsn47_1 sn47_1 sn48_1 11.551961
Rsp47_2 sp47_2 sp48_2 11.551961
Rsn47_2 sn47_2 sn48_2 11.551961
Rsp47_3 sp47_3 sp48_3 11.551961
Rsn47_3 sn47_3 sn48_3 11.551961
Rsp47_4 sp47_4 sp48_4 11.551961
Rsn47_4 sn47_4 sn48_4 11.551961
Rsp47_5 sp47_5 sp48_5 11.551961
Rsn47_5 sn47_5 sn48_5 11.551961
Rsp47_6 sp47_6 sp48_6 11.551961
Rsn47_6 sn47_6 sn48_6 11.551961
Rsp47_7 sp47_7 sp48_7 11.551961
Rsn47_7 sn47_7 sn48_7 11.551961
Rsp47_8 sp47_8 sp48_8 11.551961
Rsn47_8 sn47_8 sn48_8 11.551961
Rsp47_9 sp47_9 sp48_9 11.551961
Rsn47_9 sn47_9 sn48_9 11.551961
Rsp47_10 sp47_10 sp48_10 11.551961
Rsn47_10 sn47_10 sn48_10 11.551961
Rsp48_1 sp48_1 sp49_1 11.551961
Rsn48_1 sn48_1 sn49_1 11.551961
Rsp48_2 sp48_2 sp49_2 11.551961
Rsn48_2 sn48_2 sn49_2 11.551961
Rsp48_3 sp48_3 sp49_3 11.551961
Rsn48_3 sn48_3 sn49_3 11.551961
Rsp48_4 sp48_4 sp49_4 11.551961
Rsn48_4 sn48_4 sn49_4 11.551961
Rsp48_5 sp48_5 sp49_5 11.551961
Rsn48_5 sn48_5 sn49_5 11.551961
Rsp48_6 sp48_6 sp49_6 11.551961
Rsn48_6 sn48_6 sn49_6 11.551961
Rsp48_7 sp48_7 sp49_7 11.551961
Rsn48_7 sn48_7 sn49_7 11.551961
Rsp48_8 sp48_8 sp49_8 11.551961
Rsn48_8 sn48_8 sn49_8 11.551961
Rsp48_9 sp48_9 sp49_9 11.551961
Rsn48_9 sn48_9 sn49_9 11.551961
Rsp48_10 sp48_10 sp49_10 11.551961
Rsn48_10 sn48_10 sn49_10 11.551961
Rsp49_1 sp49_1 sp50_1 11.551961
Rsn49_1 sn49_1 sn50_1 11.551961
Rsp49_2 sp49_2 sp50_2 11.551961
Rsn49_2 sn49_2 sn50_2 11.551961
Rsp49_3 sp49_3 sp50_3 11.551961
Rsn49_3 sn49_3 sn50_3 11.551961
Rsp49_4 sp49_4 sp50_4 11.551961
Rsn49_4 sn49_4 sn50_4 11.551961
Rsp49_5 sp49_5 sp50_5 11.551961
Rsn49_5 sn49_5 sn50_5 11.551961
Rsp49_6 sp49_6 sp50_6 11.551961
Rsn49_6 sn49_6 sn50_6 11.551961
Rsp49_7 sp49_7 sp50_7 11.551961
Rsn49_7 sn49_7 sn50_7 11.551961
Rsp49_8 sp49_8 sp50_8 11.551961
Rsn49_8 sn49_8 sn50_8 11.551961
Rsp49_9 sp49_9 sp50_9 11.551961
Rsn49_9 sn49_9 sn50_9 11.551961
Rsp49_10 sp49_10 sp50_10 11.551961
Rsn49_10 sn49_10 sn50_10 11.551961
Rsp50_1 sp50_1 sp51_1 11.551961
Rsn50_1 sn50_1 sn51_1 11.551961
Rsp50_2 sp50_2 sp51_2 11.551961
Rsn50_2 sn50_2 sn51_2 11.551961
Rsp50_3 sp50_3 sp51_3 11.551961
Rsn50_3 sn50_3 sn51_3 11.551961
Rsp50_4 sp50_4 sp51_4 11.551961
Rsn50_4 sn50_4 sn51_4 11.551961
Rsp50_5 sp50_5 sp51_5 11.551961
Rsn50_5 sn50_5 sn51_5 11.551961
Rsp50_6 sp50_6 sp51_6 11.551961
Rsn50_6 sn50_6 sn51_6 11.551961
Rsp50_7 sp50_7 sp51_7 11.551961
Rsn50_7 sn50_7 sn51_7 11.551961
Rsp50_8 sp50_8 sp51_8 11.551961
Rsn50_8 sn50_8 sn51_8 11.551961
Rsp50_9 sp50_9 sp51_9 11.551961
Rsn50_9 sn50_9 sn51_9 11.551961
Rsp50_10 sp50_10 sp51_10 11.551961
Rsn50_10 sn50_10 sn51_10 11.551961
Rsp51_1 sp51_1 sp52_1 11.551961
Rsn51_1 sn51_1 sn52_1 11.551961
Rsp51_2 sp51_2 sp52_2 11.551961
Rsn51_2 sn51_2 sn52_2 11.551961
Rsp51_3 sp51_3 sp52_3 11.551961
Rsn51_3 sn51_3 sn52_3 11.551961
Rsp51_4 sp51_4 sp52_4 11.551961
Rsn51_4 sn51_4 sn52_4 11.551961
Rsp51_5 sp51_5 sp52_5 11.551961
Rsn51_5 sn51_5 sn52_5 11.551961
Rsp51_6 sp51_6 sp52_6 11.551961
Rsn51_6 sn51_6 sn52_6 11.551961
Rsp51_7 sp51_7 sp52_7 11.551961
Rsn51_7 sn51_7 sn52_7 11.551961
Rsp51_8 sp51_8 sp52_8 11.551961
Rsn51_8 sn51_8 sn52_8 11.551961
Rsp51_9 sp51_9 sp52_9 11.551961
Rsn51_9 sn51_9 sn52_9 11.551961
Rsp51_10 sp51_10 sp52_10 11.551961
Rsn51_10 sn51_10 sn52_10 11.551961
Rsp52_1 sp52_1 sp53_1 11.551961
Rsn52_1 sn52_1 sn53_1 11.551961
Rsp52_2 sp52_2 sp53_2 11.551961
Rsn52_2 sn52_2 sn53_2 11.551961
Rsp52_3 sp52_3 sp53_3 11.551961
Rsn52_3 sn52_3 sn53_3 11.551961
Rsp52_4 sp52_4 sp53_4 11.551961
Rsn52_4 sn52_4 sn53_4 11.551961
Rsp52_5 sp52_5 sp53_5 11.551961
Rsn52_5 sn52_5 sn53_5 11.551961
Rsp52_6 sp52_6 sp53_6 11.551961
Rsn52_6 sn52_6 sn53_6 11.551961
Rsp52_7 sp52_7 sp53_7 11.551961
Rsn52_7 sn52_7 sn53_7 11.551961
Rsp52_8 sp52_8 sp53_8 11.551961
Rsn52_8 sn52_8 sn53_8 11.551961
Rsp52_9 sp52_9 sp53_9 11.551961
Rsn52_9 sn52_9 sn53_9 11.551961
Rsp52_10 sp52_10 sp53_10 11.551961
Rsn52_10 sn52_10 sn53_10 11.551961
Rsp53_1 sp53_1 sp54_1 11.551961
Rsn53_1 sn53_1 sn54_1 11.551961
Rsp53_2 sp53_2 sp54_2 11.551961
Rsn53_2 sn53_2 sn54_2 11.551961
Rsp53_3 sp53_3 sp54_3 11.551961
Rsn53_3 sn53_3 sn54_3 11.551961
Rsp53_4 sp53_4 sp54_4 11.551961
Rsn53_4 sn53_4 sn54_4 11.551961
Rsp53_5 sp53_5 sp54_5 11.551961
Rsn53_5 sn53_5 sn54_5 11.551961
Rsp53_6 sp53_6 sp54_6 11.551961
Rsn53_6 sn53_6 sn54_6 11.551961
Rsp53_7 sp53_7 sp54_7 11.551961
Rsn53_7 sn53_7 sn54_7 11.551961
Rsp53_8 sp53_8 sp54_8 11.551961
Rsn53_8 sn53_8 sn54_8 11.551961
Rsp53_9 sp53_9 sp54_9 11.551961
Rsn53_9 sn53_9 sn54_9 11.551961
Rsp53_10 sp53_10 sp54_10 11.551961
Rsn53_10 sn53_10 sn54_10 11.551961
Rsp54_1 sp54_1 sp55_1 11.551961
Rsn54_1 sn54_1 sn55_1 11.551961
Rsp54_2 sp54_2 sp55_2 11.551961
Rsn54_2 sn54_2 sn55_2 11.551961
Rsp54_3 sp54_3 sp55_3 11.551961
Rsn54_3 sn54_3 sn55_3 11.551961
Rsp54_4 sp54_4 sp55_4 11.551961
Rsn54_4 sn54_4 sn55_4 11.551961
Rsp54_5 sp54_5 sp55_5 11.551961
Rsn54_5 sn54_5 sn55_5 11.551961
Rsp54_6 sp54_6 sp55_6 11.551961
Rsn54_6 sn54_6 sn55_6 11.551961
Rsp54_7 sp54_7 sp55_7 11.551961
Rsn54_7 sn54_7 sn55_7 11.551961
Rsp54_8 sp54_8 sp55_8 11.551961
Rsn54_8 sn54_8 sn55_8 11.551961
Rsp54_9 sp54_9 sp55_9 11.551961
Rsn54_9 sn54_9 sn55_9 11.551961
Rsp54_10 sp54_10 sp55_10 11.551961
Rsn54_10 sn54_10 sn55_10 11.551961
Rsp55_1 sp55_1 sp56_1 11.551961
Rsn55_1 sn55_1 sn56_1 11.551961
Rsp55_2 sp55_2 sp56_2 11.551961
Rsn55_2 sn55_2 sn56_2 11.551961
Rsp55_3 sp55_3 sp56_3 11.551961
Rsn55_3 sn55_3 sn56_3 11.551961
Rsp55_4 sp55_4 sp56_4 11.551961
Rsn55_4 sn55_4 sn56_4 11.551961
Rsp55_5 sp55_5 sp56_5 11.551961
Rsn55_5 sn55_5 sn56_5 11.551961
Rsp55_6 sp55_6 sp56_6 11.551961
Rsn55_6 sn55_6 sn56_6 11.551961
Rsp55_7 sp55_7 sp56_7 11.551961
Rsn55_7 sn55_7 sn56_7 11.551961
Rsp55_8 sp55_8 sp56_8 11.551961
Rsn55_8 sn55_8 sn56_8 11.551961
Rsp55_9 sp55_9 sp56_9 11.551961
Rsn55_9 sn55_9 sn56_9 11.551961
Rsp55_10 sp55_10 sp56_10 11.551961
Rsn55_10 sn55_10 sn56_10 11.551961
Rsp56_1 sp56_1 sp57_1 11.551961
Rsn56_1 sn56_1 sn57_1 11.551961
Rsp56_2 sp56_2 sp57_2 11.551961
Rsn56_2 sn56_2 sn57_2 11.551961
Rsp56_3 sp56_3 sp57_3 11.551961
Rsn56_3 sn56_3 sn57_3 11.551961
Rsp56_4 sp56_4 sp57_4 11.551961
Rsn56_4 sn56_4 sn57_4 11.551961
Rsp56_5 sp56_5 sp57_5 11.551961
Rsn56_5 sn56_5 sn57_5 11.551961
Rsp56_6 sp56_6 sp57_6 11.551961
Rsn56_6 sn56_6 sn57_6 11.551961
Rsp56_7 sp56_7 sp57_7 11.551961
Rsn56_7 sn56_7 sn57_7 11.551961
Rsp56_8 sp56_8 sp57_8 11.551961
Rsn56_8 sn56_8 sn57_8 11.551961
Rsp56_9 sp56_9 sp57_9 11.551961
Rsn56_9 sn56_9 sn57_9 11.551961
Rsp56_10 sp56_10 sp57_10 11.551961
Rsn56_10 sn56_10 sn57_10 11.551961
Rsp57_1 sp57_1 sp1_p2 11.551961
Rsn57_1 sn57_1 sn1_p2 11.551961
Rsp57_2 sp57_2 sp2_p2 11.551961
Rsn57_2 sn57_2 sn2_p2 11.551961
Rsp57_3 sp57_3 sp3_p2 11.551961
Rsn57_3 sn57_3 sn3_p2 11.551961
Rsp57_4 sp57_4 sp4_p2 11.551961
Rsn57_4 sn57_4 sn4_p2 11.551961
Rsp57_5 sp57_5 sp5_p2 11.551961
Rsn57_5 sn57_5 sn5_p2 11.551961
Rsp57_6 sp57_6 sp6_p2 11.551961
Rsn57_6 sn57_6 sn6_p2 11.551961
Rsp57_7 sp57_7 sp7_p2 11.551961
Rsn57_7 sn57_7 sn7_p2 11.551961
Rsp57_8 sp57_8 sp8_p2 11.551961
Rsn57_8 sn57_8 sn8_p2 11.551961
Rsp57_9 sp57_9 sp9_p2 11.551961
Rsn57_9 sn57_9 sn9_p2 11.551961
Rsp57_10 sp57_10 sp10_p2 11.551961
Rsn57_10 sn57_10 sn10_p2 11.551961
Rsp58_1 sp58_1 sp59_1 11.551961
Rsn58_1 sn58_1 sn59_1 11.551961
Rsp58_2 sp58_2 sp59_2 11.551961
Rsn58_2 sn58_2 sn59_2 11.551961
Rsp58_3 sp58_3 sp59_3 11.551961
Rsn58_3 sn58_3 sn59_3 11.551961
Rsp58_4 sp58_4 sp59_4 11.551961
Rsn58_4 sn58_4 sn59_4 11.551961
Rsp58_5 sp58_5 sp59_5 11.551961
Rsn58_5 sn58_5 sn59_5 11.551961
Rsp58_6 sp58_6 sp59_6 11.551961
Rsn58_6 sn58_6 sn59_6 11.551961
Rsp58_7 sp58_7 sp59_7 11.551961
Rsn58_7 sn58_7 sn59_7 11.551961
Rsp58_8 sp58_8 sp59_8 11.551961
Rsn58_8 sn58_8 sn59_8 11.551961
Rsp58_9 sp58_9 sp59_9 11.551961
Rsn58_9 sn58_9 sn59_9 11.551961
Rsp58_10 sp58_10 sp59_10 11.551961
Rsn58_10 sn58_10 sn59_10 11.551961
Rsp59_1 sp59_1 sp60_1 11.551961
Rsn59_1 sn59_1 sn60_1 11.551961
Rsp59_2 sp59_2 sp60_2 11.551961
Rsn59_2 sn59_2 sn60_2 11.551961
Rsp59_3 sp59_3 sp60_3 11.551961
Rsn59_3 sn59_3 sn60_3 11.551961
Rsp59_4 sp59_4 sp60_4 11.551961
Rsn59_4 sn59_4 sn60_4 11.551961
Rsp59_5 sp59_5 sp60_5 11.551961
Rsn59_5 sn59_5 sn60_5 11.551961
Rsp59_6 sp59_6 sp60_6 11.551961
Rsn59_6 sn59_6 sn60_6 11.551961
Rsp59_7 sp59_7 sp60_7 11.551961
Rsn59_7 sn59_7 sn60_7 11.551961
Rsp59_8 sp59_8 sp60_8 11.551961
Rsn59_8 sn59_8 sn60_8 11.551961
Rsp59_9 sp59_9 sp60_9 11.551961
Rsn59_9 sn59_9 sn60_9 11.551961
Rsp59_10 sp59_10 sp60_10 11.551961
Rsn59_10 sn59_10 sn60_10 11.551961
Rsp60_1 sp60_1 sp61_1 11.551961
Rsn60_1 sn60_1 sn61_1 11.551961
Rsp60_2 sp60_2 sp61_2 11.551961
Rsn60_2 sn60_2 sn61_2 11.551961
Rsp60_3 sp60_3 sp61_3 11.551961
Rsn60_3 sn60_3 sn61_3 11.551961
Rsp60_4 sp60_4 sp61_4 11.551961
Rsn60_4 sn60_4 sn61_4 11.551961
Rsp60_5 sp60_5 sp61_5 11.551961
Rsn60_5 sn60_5 sn61_5 11.551961
Rsp60_6 sp60_6 sp61_6 11.551961
Rsn60_6 sn60_6 sn61_6 11.551961
Rsp60_7 sp60_7 sp61_7 11.551961
Rsn60_7 sn60_7 sn61_7 11.551961
Rsp60_8 sp60_8 sp61_8 11.551961
Rsn60_8 sn60_8 sn61_8 11.551961
Rsp60_9 sp60_9 sp61_9 11.551961
Rsn60_9 sn60_9 sn61_9 11.551961
Rsp60_10 sp60_10 sp61_10 11.551961
Rsn60_10 sn60_10 sn61_10 11.551961
Rsp61_1 sp61_1 sp62_1 11.551961
Rsn61_1 sn61_1 sn62_1 11.551961
Rsp61_2 sp61_2 sp62_2 11.551961
Rsn61_2 sn61_2 sn62_2 11.551961
Rsp61_3 sp61_3 sp62_3 11.551961
Rsn61_3 sn61_3 sn62_3 11.551961
Rsp61_4 sp61_4 sp62_4 11.551961
Rsn61_4 sn61_4 sn62_4 11.551961
Rsp61_5 sp61_5 sp62_5 11.551961
Rsn61_5 sn61_5 sn62_5 11.551961
Rsp61_6 sp61_6 sp62_6 11.551961
Rsn61_6 sn61_6 sn62_6 11.551961
Rsp61_7 sp61_7 sp62_7 11.551961
Rsn61_7 sn61_7 sn62_7 11.551961
Rsp61_8 sp61_8 sp62_8 11.551961
Rsn61_8 sn61_8 sn62_8 11.551961
Rsp61_9 sp61_9 sp62_9 11.551961
Rsn61_9 sn61_9 sn62_9 11.551961
Rsp61_10 sp61_10 sp62_10 11.551961
Rsn61_10 sn61_10 sn62_10 11.551961
Rsp62_1 sp62_1 sp63_1 11.551961
Rsn62_1 sn62_1 sn63_1 11.551961
Rsp62_2 sp62_2 sp63_2 11.551961
Rsn62_2 sn62_2 sn63_2 11.551961
Rsp62_3 sp62_3 sp63_3 11.551961
Rsn62_3 sn62_3 sn63_3 11.551961
Rsp62_4 sp62_4 sp63_4 11.551961
Rsn62_4 sn62_4 sn63_4 11.551961
Rsp62_5 sp62_5 sp63_5 11.551961
Rsn62_5 sn62_5 sn63_5 11.551961
Rsp62_6 sp62_6 sp63_6 11.551961
Rsn62_6 sn62_6 sn63_6 11.551961
Rsp62_7 sp62_7 sp63_7 11.551961
Rsn62_7 sn62_7 sn63_7 11.551961
Rsp62_8 sp62_8 sp63_8 11.551961
Rsn62_8 sn62_8 sn63_8 11.551961
Rsp62_9 sp62_9 sp63_9 11.551961
Rsn62_9 sn62_9 sn63_9 11.551961
Rsp62_10 sp62_10 sp63_10 11.551961
Rsn62_10 sn62_10 sn63_10 11.551961
Rsp63_1 sp63_1 sp64_1 11.551961
Rsn63_1 sn63_1 sn64_1 11.551961
Rsp63_2 sp63_2 sp64_2 11.551961
Rsn63_2 sn63_2 sn64_2 11.551961
Rsp63_3 sp63_3 sp64_3 11.551961
Rsn63_3 sn63_3 sn64_3 11.551961
Rsp63_4 sp63_4 sp64_4 11.551961
Rsn63_4 sn63_4 sn64_4 11.551961
Rsp63_5 sp63_5 sp64_5 11.551961
Rsn63_5 sn63_5 sn64_5 11.551961
Rsp63_6 sp63_6 sp64_6 11.551961
Rsn63_6 sn63_6 sn64_6 11.551961
Rsp63_7 sp63_7 sp64_7 11.551961
Rsn63_7 sn63_7 sn64_7 11.551961
Rsp63_8 sp63_8 sp64_8 11.551961
Rsn63_8 sn63_8 sn64_8 11.551961
Rsp63_9 sp63_9 sp64_9 11.551961
Rsn63_9 sn63_9 sn64_9 11.551961
Rsp63_10 sp63_10 sp64_10 11.551961
Rsn63_10 sn63_10 sn64_10 11.551961
Rsp64_1 sp64_1 sp65_1 11.551961
Rsn64_1 sn64_1 sn65_1 11.551961
Rsp64_2 sp64_2 sp65_2 11.551961
Rsn64_2 sn64_2 sn65_2 11.551961
Rsp64_3 sp64_3 sp65_3 11.551961
Rsn64_3 sn64_3 sn65_3 11.551961
Rsp64_4 sp64_4 sp65_4 11.551961
Rsn64_4 sn64_4 sn65_4 11.551961
Rsp64_5 sp64_5 sp65_5 11.551961
Rsn64_5 sn64_5 sn65_5 11.551961
Rsp64_6 sp64_6 sp65_6 11.551961
Rsn64_6 sn64_6 sn65_6 11.551961
Rsp64_7 sp64_7 sp65_7 11.551961
Rsn64_7 sn64_7 sn65_7 11.551961
Rsp64_8 sp64_8 sp65_8 11.551961
Rsn64_8 sn64_8 sn65_8 11.551961
Rsp64_9 sp64_9 sp65_9 11.551961
Rsn64_9 sn64_9 sn65_9 11.551961
Rsp64_10 sp64_10 sp65_10 11.551961
Rsn64_10 sn64_10 sn65_10 11.551961
Rsp65_1 sp65_1 sp66_1 11.551961
Rsn65_1 sn65_1 sn66_1 11.551961
Rsp65_2 sp65_2 sp66_2 11.551961
Rsn65_2 sn65_2 sn66_2 11.551961
Rsp65_3 sp65_3 sp66_3 11.551961
Rsn65_3 sn65_3 sn66_3 11.551961
Rsp65_4 sp65_4 sp66_4 11.551961
Rsn65_4 sn65_4 sn66_4 11.551961
Rsp65_5 sp65_5 sp66_5 11.551961
Rsn65_5 sn65_5 sn66_5 11.551961
Rsp65_6 sp65_6 sp66_6 11.551961
Rsn65_6 sn65_6 sn66_6 11.551961
Rsp65_7 sp65_7 sp66_7 11.551961
Rsn65_7 sn65_7 sn66_7 11.551961
Rsp65_8 sp65_8 sp66_8 11.551961
Rsn65_8 sn65_8 sn66_8 11.551961
Rsp65_9 sp65_9 sp66_9 11.551961
Rsn65_9 sn65_9 sn66_9 11.551961
Rsp65_10 sp65_10 sp66_10 11.551961
Rsn65_10 sn65_10 sn66_10 11.551961
Rsp66_1 sp66_1 sp67_1 11.551961
Rsn66_1 sn66_1 sn67_1 11.551961
Rsp66_2 sp66_2 sp67_2 11.551961
Rsn66_2 sn66_2 sn67_2 11.551961
Rsp66_3 sp66_3 sp67_3 11.551961
Rsn66_3 sn66_3 sn67_3 11.551961
Rsp66_4 sp66_4 sp67_4 11.551961
Rsn66_4 sn66_4 sn67_4 11.551961
Rsp66_5 sp66_5 sp67_5 11.551961
Rsn66_5 sn66_5 sn67_5 11.551961
Rsp66_6 sp66_6 sp67_6 11.551961
Rsn66_6 sn66_6 sn67_6 11.551961
Rsp66_7 sp66_7 sp67_7 11.551961
Rsn66_7 sn66_7 sn67_7 11.551961
Rsp66_8 sp66_8 sp67_8 11.551961
Rsn66_8 sn66_8 sn67_8 11.551961
Rsp66_9 sp66_9 sp67_9 11.551961
Rsn66_9 sn66_9 sn67_9 11.551961
Rsp66_10 sp66_10 sp67_10 11.551961
Rsn66_10 sn66_10 sn67_10 11.551961
Rsp67_1 sp67_1 sp68_1 11.551961
Rsn67_1 sn67_1 sn68_1 11.551961
Rsp67_2 sp67_2 sp68_2 11.551961
Rsn67_2 sn67_2 sn68_2 11.551961
Rsp67_3 sp67_3 sp68_3 11.551961
Rsn67_3 sn67_3 sn68_3 11.551961
Rsp67_4 sp67_4 sp68_4 11.551961
Rsn67_4 sn67_4 sn68_4 11.551961
Rsp67_5 sp67_5 sp68_5 11.551961
Rsn67_5 sn67_5 sn68_5 11.551961
Rsp67_6 sp67_6 sp68_6 11.551961
Rsn67_6 sn67_6 sn68_6 11.551961
Rsp67_7 sp67_7 sp68_7 11.551961
Rsn67_7 sn67_7 sn68_7 11.551961
Rsp67_8 sp67_8 sp68_8 11.551961
Rsn67_8 sn67_8 sn68_8 11.551961
Rsp67_9 sp67_9 sp68_9 11.551961
Rsn67_9 sn67_9 sn68_9 11.551961
Rsp67_10 sp67_10 sp68_10 11.551961
Rsn67_10 sn67_10 sn68_10 11.551961
Rsp68_1 sp68_1 sp69_1 11.551961
Rsn68_1 sn68_1 sn69_1 11.551961
Rsp68_2 sp68_2 sp69_2 11.551961
Rsn68_2 sn68_2 sn69_2 11.551961
Rsp68_3 sp68_3 sp69_3 11.551961
Rsn68_3 sn68_3 sn69_3 11.551961
Rsp68_4 sp68_4 sp69_4 11.551961
Rsn68_4 sn68_4 sn69_4 11.551961
Rsp68_5 sp68_5 sp69_5 11.551961
Rsn68_5 sn68_5 sn69_5 11.551961
Rsp68_6 sp68_6 sp69_6 11.551961
Rsn68_6 sn68_6 sn69_6 11.551961
Rsp68_7 sp68_7 sp69_7 11.551961
Rsn68_7 sn68_7 sn69_7 11.551961
Rsp68_8 sp68_8 sp69_8 11.551961
Rsn68_8 sn68_8 sn69_8 11.551961
Rsp68_9 sp68_9 sp69_9 11.551961
Rsn68_9 sn68_9 sn69_9 11.551961
Rsp68_10 sp68_10 sp69_10 11.551961
Rsn68_10 sn68_10 sn69_10 11.551961
Rsp69_1 sp69_1 sp70_1 11.551961
Rsn69_1 sn69_1 sn70_1 11.551961
Rsp69_2 sp69_2 sp70_2 11.551961
Rsn69_2 sn69_2 sn70_2 11.551961
Rsp69_3 sp69_3 sp70_3 11.551961
Rsn69_3 sn69_3 sn70_3 11.551961
Rsp69_4 sp69_4 sp70_4 11.551961
Rsn69_4 sn69_4 sn70_4 11.551961
Rsp69_5 sp69_5 sp70_5 11.551961
Rsn69_5 sn69_5 sn70_5 11.551961
Rsp69_6 sp69_6 sp70_6 11.551961
Rsn69_6 sn69_6 sn70_6 11.551961
Rsp69_7 sp69_7 sp70_7 11.551961
Rsn69_7 sn69_7 sn70_7 11.551961
Rsp69_8 sp69_8 sp70_8 11.551961
Rsn69_8 sn69_8 sn70_8 11.551961
Rsp69_9 sp69_9 sp70_9 11.551961
Rsn69_9 sn69_9 sn70_9 11.551961
Rsp69_10 sp69_10 sp70_10 11.551961
Rsn69_10 sn69_10 sn70_10 11.551961
Rsp70_1 sp70_1 sp71_1 11.551961
Rsn70_1 sn70_1 sn71_1 11.551961
Rsp70_2 sp70_2 sp71_2 11.551961
Rsn70_2 sn70_2 sn71_2 11.551961
Rsp70_3 sp70_3 sp71_3 11.551961
Rsn70_3 sn70_3 sn71_3 11.551961
Rsp70_4 sp70_4 sp71_4 11.551961
Rsn70_4 sn70_4 sn71_4 11.551961
Rsp70_5 sp70_5 sp71_5 11.551961
Rsn70_5 sn70_5 sn71_5 11.551961
Rsp70_6 sp70_6 sp71_6 11.551961
Rsn70_6 sn70_6 sn71_6 11.551961
Rsp70_7 sp70_7 sp71_7 11.551961
Rsn70_7 sn70_7 sn71_7 11.551961
Rsp70_8 sp70_8 sp71_8 11.551961
Rsn70_8 sn70_8 sn71_8 11.551961
Rsp70_9 sp70_9 sp71_9 11.551961
Rsn70_9 sn70_9 sn71_9 11.551961
Rsp70_10 sp70_10 sp71_10 11.551961
Rsn70_10 sn70_10 sn71_10 11.551961
Rsp71_1 sp71_1 sp72_1 11.551961
Rsn71_1 sn71_1 sn72_1 11.551961
Rsp71_2 sp71_2 sp72_2 11.551961
Rsn71_2 sn71_2 sn72_2 11.551961
Rsp71_3 sp71_3 sp72_3 11.551961
Rsn71_3 sn71_3 sn72_3 11.551961
Rsp71_4 sp71_4 sp72_4 11.551961
Rsn71_4 sn71_4 sn72_4 11.551961
Rsp71_5 sp71_5 sp72_5 11.551961
Rsn71_5 sn71_5 sn72_5 11.551961
Rsp71_6 sp71_6 sp72_6 11.551961
Rsn71_6 sn71_6 sn72_6 11.551961
Rsp71_7 sp71_7 sp72_7 11.551961
Rsn71_7 sn71_7 sn72_7 11.551961
Rsp71_8 sp71_8 sp72_8 11.551961
Rsn71_8 sn71_8 sn72_8 11.551961
Rsp71_9 sp71_9 sp72_9 11.551961
Rsn71_9 sn71_9 sn72_9 11.551961
Rsp71_10 sp71_10 sp72_10 11.551961
Rsn71_10 sn71_10 sn72_10 11.551961
Rsp72_1 sp72_1 sp73_1 11.551961
Rsn72_1 sn72_1 sn73_1 11.551961
Rsp72_2 sp72_2 sp73_2 11.551961
Rsn72_2 sn72_2 sn73_2 11.551961
Rsp72_3 sp72_3 sp73_3 11.551961
Rsn72_3 sn72_3 sn73_3 11.551961
Rsp72_4 sp72_4 sp73_4 11.551961
Rsn72_4 sn72_4 sn73_4 11.551961
Rsp72_5 sp72_5 sp73_5 11.551961
Rsn72_5 sn72_5 sn73_5 11.551961
Rsp72_6 sp72_6 sp73_6 11.551961
Rsn72_6 sn72_6 sn73_6 11.551961
Rsp72_7 sp72_7 sp73_7 11.551961
Rsn72_7 sn72_7 sn73_7 11.551961
Rsp72_8 sp72_8 sp73_8 11.551961
Rsn72_8 sn72_8 sn73_8 11.551961
Rsp72_9 sp72_9 sp73_9 11.551961
Rsn72_9 sn72_9 sn73_9 11.551961
Rsp72_10 sp72_10 sp73_10 11.551961
Rsn72_10 sn72_10 sn73_10 11.551961
Rsp73_1 sp73_1 sp74_1 11.551961
Rsn73_1 sn73_1 sn74_1 11.551961
Rsp73_2 sp73_2 sp74_2 11.551961
Rsn73_2 sn73_2 sn74_2 11.551961
Rsp73_3 sp73_3 sp74_3 11.551961
Rsn73_3 sn73_3 sn74_3 11.551961
Rsp73_4 sp73_4 sp74_4 11.551961
Rsn73_4 sn73_4 sn74_4 11.551961
Rsp73_5 sp73_5 sp74_5 11.551961
Rsn73_5 sn73_5 sn74_5 11.551961
Rsp73_6 sp73_6 sp74_6 11.551961
Rsn73_6 sn73_6 sn74_6 11.551961
Rsp73_7 sp73_7 sp74_7 11.551961
Rsn73_7 sn73_7 sn74_7 11.551961
Rsp73_8 sp73_8 sp74_8 11.551961
Rsn73_8 sn73_8 sn74_8 11.551961
Rsp73_9 sp73_9 sp74_9 11.551961
Rsn73_9 sn73_9 sn74_9 11.551961
Rsp73_10 sp73_10 sp74_10 11.551961
Rsn73_10 sn73_10 sn74_10 11.551961
Rsp74_1 sp74_1 sp75_1 11.551961
Rsn74_1 sn74_1 sn75_1 11.551961
Rsp74_2 sp74_2 sp75_2 11.551961
Rsn74_2 sn74_2 sn75_2 11.551961
Rsp74_3 sp74_3 sp75_3 11.551961
Rsn74_3 sn74_3 sn75_3 11.551961
Rsp74_4 sp74_4 sp75_4 11.551961
Rsn74_4 sn74_4 sn75_4 11.551961
Rsp74_5 sp74_5 sp75_5 11.551961
Rsn74_5 sn74_5 sn75_5 11.551961
Rsp74_6 sp74_6 sp75_6 11.551961
Rsn74_6 sn74_6 sn75_6 11.551961
Rsp74_7 sp74_7 sp75_7 11.551961
Rsn74_7 sn74_7 sn75_7 11.551961
Rsp74_8 sp74_8 sp75_8 11.551961
Rsn74_8 sn74_8 sn75_8 11.551961
Rsp74_9 sp74_9 sp75_9 11.551961
Rsn74_9 sn74_9 sn75_9 11.551961
Rsp74_10 sp74_10 sp75_10 11.551961
Rsn74_10 sn74_10 sn75_10 11.551961
Rsp75_1 sp75_1 sp76_1 11.551961
Rsn75_1 sn75_1 sn76_1 11.551961
Rsp75_2 sp75_2 sp76_2 11.551961
Rsn75_2 sn75_2 sn76_2 11.551961
Rsp75_3 sp75_3 sp76_3 11.551961
Rsn75_3 sn75_3 sn76_3 11.551961
Rsp75_4 sp75_4 sp76_4 11.551961
Rsn75_4 sn75_4 sn76_4 11.551961
Rsp75_5 sp75_5 sp76_5 11.551961
Rsn75_5 sn75_5 sn76_5 11.551961
Rsp75_6 sp75_6 sp76_6 11.551961
Rsn75_6 sn75_6 sn76_6 11.551961
Rsp75_7 sp75_7 sp76_7 11.551961
Rsn75_7 sn75_7 sn76_7 11.551961
Rsp75_8 sp75_8 sp76_8 11.551961
Rsn75_8 sn75_8 sn76_8 11.551961
Rsp75_9 sp75_9 sp76_9 11.551961
Rsn75_9 sn75_9 sn76_9 11.551961
Rsp75_10 sp75_10 sp76_10 11.551961
Rsn75_10 sn75_10 sn76_10 11.551961
Rsp76_1 sp76_1 sp77_1 11.551961
Rsn76_1 sn76_1 sn77_1 11.551961
Rsp76_2 sp76_2 sp77_2 11.551961
Rsn76_2 sn76_2 sn77_2 11.551961
Rsp76_3 sp76_3 sp77_3 11.551961
Rsn76_3 sn76_3 sn77_3 11.551961
Rsp76_4 sp76_4 sp77_4 11.551961
Rsn76_4 sn76_4 sn77_4 11.551961
Rsp76_5 sp76_5 sp77_5 11.551961
Rsn76_5 sn76_5 sn77_5 11.551961
Rsp76_6 sp76_6 sp77_6 11.551961
Rsn76_6 sn76_6 sn77_6 11.551961
Rsp76_7 sp76_7 sp77_7 11.551961
Rsn76_7 sn76_7 sn77_7 11.551961
Rsp76_8 sp76_8 sp77_8 11.551961
Rsn76_8 sn76_8 sn77_8 11.551961
Rsp76_9 sp76_9 sp77_9 11.551961
Rsn76_9 sn76_9 sn77_9 11.551961
Rsp76_10 sp76_10 sp77_10 11.551961
Rsn76_10 sn76_10 sn77_10 11.551961
Rsp77_1 sp77_1 sp78_1 11.551961
Rsn77_1 sn77_1 sn78_1 11.551961
Rsp77_2 sp77_2 sp78_2 11.551961
Rsn77_2 sn77_2 sn78_2 11.551961
Rsp77_3 sp77_3 sp78_3 11.551961
Rsn77_3 sn77_3 sn78_3 11.551961
Rsp77_4 sp77_4 sp78_4 11.551961
Rsn77_4 sn77_4 sn78_4 11.551961
Rsp77_5 sp77_5 sp78_5 11.551961
Rsn77_5 sn77_5 sn78_5 11.551961
Rsp77_6 sp77_6 sp78_6 11.551961
Rsn77_6 sn77_6 sn78_6 11.551961
Rsp77_7 sp77_7 sp78_7 11.551961
Rsn77_7 sn77_7 sn78_7 11.551961
Rsp77_8 sp77_8 sp78_8 11.551961
Rsn77_8 sn77_8 sn78_8 11.551961
Rsp77_9 sp77_9 sp78_9 11.551961
Rsn77_9 sn77_9 sn78_9 11.551961
Rsp77_10 sp77_10 sp78_10 11.551961
Rsn77_10 sn77_10 sn78_10 11.551961
Rsp78_1 sp78_1 sp79_1 11.551961
Rsn78_1 sn78_1 sn79_1 11.551961
Rsp78_2 sp78_2 sp79_2 11.551961
Rsn78_2 sn78_2 sn79_2 11.551961
Rsp78_3 sp78_3 sp79_3 11.551961
Rsn78_3 sn78_3 sn79_3 11.551961
Rsp78_4 sp78_4 sp79_4 11.551961
Rsn78_4 sn78_4 sn79_4 11.551961
Rsp78_5 sp78_5 sp79_5 11.551961
Rsn78_5 sn78_5 sn79_5 11.551961
Rsp78_6 sp78_6 sp79_6 11.551961
Rsn78_6 sn78_6 sn79_6 11.551961
Rsp78_7 sp78_7 sp79_7 11.551961
Rsn78_7 sn78_7 sn79_7 11.551961
Rsp78_8 sp78_8 sp79_8 11.551961
Rsn78_8 sn78_8 sn79_8 11.551961
Rsp78_9 sp78_9 sp79_9 11.551961
Rsn78_9 sn78_9 sn79_9 11.551961
Rsp78_10 sp78_10 sp79_10 11.551961
Rsn78_10 sn78_10 sn79_10 11.551961
Rsp79_1 sp79_1 sp80_1 11.551961
Rsn79_1 sn79_1 sn80_1 11.551961
Rsp79_2 sp79_2 sp80_2 11.551961
Rsn79_2 sn79_2 sn80_2 11.551961
Rsp79_3 sp79_3 sp80_3 11.551961
Rsn79_3 sn79_3 sn80_3 11.551961
Rsp79_4 sp79_4 sp80_4 11.551961
Rsn79_4 sn79_4 sn80_4 11.551961
Rsp79_5 sp79_5 sp80_5 11.551961
Rsn79_5 sn79_5 sn80_5 11.551961
Rsp79_6 sp79_6 sp80_6 11.551961
Rsn79_6 sn79_6 sn80_6 11.551961
Rsp79_7 sp79_7 sp80_7 11.551961
Rsn79_7 sn79_7 sn80_7 11.551961
Rsp79_8 sp79_8 sp80_8 11.551961
Rsn79_8 sn79_8 sn80_8 11.551961
Rsp79_9 sp79_9 sp80_9 11.551961
Rsn79_9 sn79_9 sn80_9 11.551961
Rsp79_10 sp79_10 sp80_10 11.551961
Rsn79_10 sn79_10 sn80_10 11.551961
Rsp80_1 sp80_1 sp81_1 11.551961
Rsn80_1 sn80_1 sn81_1 11.551961
Rsp80_2 sp80_2 sp81_2 11.551961
Rsn80_2 sn80_2 sn81_2 11.551961
Rsp80_3 sp80_3 sp81_3 11.551961
Rsn80_3 sn80_3 sn81_3 11.551961
Rsp80_4 sp80_4 sp81_4 11.551961
Rsn80_4 sn80_4 sn81_4 11.551961
Rsp80_5 sp80_5 sp81_5 11.551961
Rsn80_5 sn80_5 sn81_5 11.551961
Rsp80_6 sp80_6 sp81_6 11.551961
Rsn80_6 sn80_6 sn81_6 11.551961
Rsp80_7 sp80_7 sp81_7 11.551961
Rsn80_7 sn80_7 sn81_7 11.551961
Rsp80_8 sp80_8 sp81_8 11.551961
Rsn80_8 sn80_8 sn81_8 11.551961
Rsp80_9 sp80_9 sp81_9 11.551961
Rsn80_9 sn80_9 sn81_9 11.551961
Rsp80_10 sp80_10 sp81_10 11.551961
Rsn80_10 sn80_10 sn81_10 11.551961
Rsp81_1 sp81_1 sp82_1 11.551961
Rsn81_1 sn81_1 sn82_1 11.551961
Rsp81_2 sp81_2 sp82_2 11.551961
Rsn81_2 sn81_2 sn82_2 11.551961
Rsp81_3 sp81_3 sp82_3 11.551961
Rsn81_3 sn81_3 sn82_3 11.551961
Rsp81_4 sp81_4 sp82_4 11.551961
Rsn81_4 sn81_4 sn82_4 11.551961
Rsp81_5 sp81_5 sp82_5 11.551961
Rsn81_5 sn81_5 sn82_5 11.551961
Rsp81_6 sp81_6 sp82_6 11.551961
Rsn81_6 sn81_6 sn82_6 11.551961
Rsp81_7 sp81_7 sp82_7 11.551961
Rsn81_7 sn81_7 sn82_7 11.551961
Rsp81_8 sp81_8 sp82_8 11.551961
Rsn81_8 sn81_8 sn82_8 11.551961
Rsp81_9 sp81_9 sp82_9 11.551961
Rsn81_9 sn81_9 sn82_9 11.551961
Rsp81_10 sp81_10 sp82_10 11.551961
Rsn81_10 sn81_10 sn82_10 11.551961
Rsp82_1 sp82_1 sp83_1 11.551961
Rsn82_1 sn82_1 sn83_1 11.551961
Rsp82_2 sp82_2 sp83_2 11.551961
Rsn82_2 sn82_2 sn83_2 11.551961
Rsp82_3 sp82_3 sp83_3 11.551961
Rsn82_3 sn82_3 sn83_3 11.551961
Rsp82_4 sp82_4 sp83_4 11.551961
Rsn82_4 sn82_4 sn83_4 11.551961
Rsp82_5 sp82_5 sp83_5 11.551961
Rsn82_5 sn82_5 sn83_5 11.551961
Rsp82_6 sp82_6 sp83_6 11.551961
Rsn82_6 sn82_6 sn83_6 11.551961
Rsp82_7 sp82_7 sp83_7 11.551961
Rsn82_7 sn82_7 sn83_7 11.551961
Rsp82_8 sp82_8 sp83_8 11.551961
Rsn82_8 sn82_8 sn83_8 11.551961
Rsp82_9 sp82_9 sp83_9 11.551961
Rsn82_9 sn82_9 sn83_9 11.551961
Rsp82_10 sp82_10 sp83_10 11.551961
Rsn82_10 sn82_10 sn83_10 11.551961
Rsp83_1 sp83_1 sp84_1 11.551961
Rsn83_1 sn83_1 sn84_1 11.551961
Rsp83_2 sp83_2 sp84_2 11.551961
Rsn83_2 sn83_2 sn84_2 11.551961
Rsp83_3 sp83_3 sp84_3 11.551961
Rsn83_3 sn83_3 sn84_3 11.551961
Rsp83_4 sp83_4 sp84_4 11.551961
Rsn83_4 sn83_4 sn84_4 11.551961
Rsp83_5 sp83_5 sp84_5 11.551961
Rsn83_5 sn83_5 sn84_5 11.551961
Rsp83_6 sp83_6 sp84_6 11.551961
Rsn83_6 sn83_6 sn84_6 11.551961
Rsp83_7 sp83_7 sp84_7 11.551961
Rsn83_7 sn83_7 sn84_7 11.551961
Rsp83_8 sp83_8 sp84_8 11.551961
Rsn83_8 sn83_8 sn84_8 11.551961
Rsp83_9 sp83_9 sp84_9 11.551961
Rsn83_9 sn83_9 sn84_9 11.551961
Rsp83_10 sp83_10 sp84_10 11.551961
Rsn83_10 sn83_10 sn84_10 11.551961
Rsp84_1 sp84_1 sp85_1 11.551961
Rsn84_1 sn84_1 sn85_1 11.551961
Rsp84_2 sp84_2 sp85_2 11.551961
Rsn84_2 sn84_2 sn85_2 11.551961
Rsp84_3 sp84_3 sp85_3 11.551961
Rsn84_3 sn84_3 sn85_3 11.551961
Rsp84_4 sp84_4 sp85_4 11.551961
Rsn84_4 sn84_4 sn85_4 11.551961
Rsp84_5 sp84_5 sp85_5 11.551961
Rsn84_5 sn84_5 sn85_5 11.551961
Rsp84_6 sp84_6 sp85_6 11.551961
Rsn84_6 sn84_6 sn85_6 11.551961
Rsp84_7 sp84_7 sp85_7 11.551961
Rsn84_7 sn84_7 sn85_7 11.551961
Rsp84_8 sp84_8 sp85_8 11.551961
Rsn84_8 sn84_8 sn85_8 11.551961
Rsp84_9 sp84_9 sp85_9 11.551961
Rsn84_9 sn84_9 sn85_9 11.551961
Rsp84_10 sp84_10 sp85_10 11.551961
Rsn84_10 sn84_10 sn85_10 11.551961
Rsp85_1 sp85_1 sp1_p3 11.551961
Rsn85_1 sn85_1 sn1_p3 11.551961
Rsp85_2 sp85_2 sp2_p3 11.551961
Rsn85_2 sn85_2 sn2_p3 11.551961
Rsp85_3 sp85_3 sp3_p3 11.551961
Rsn85_3 sn85_3 sn3_p3 11.551961
Rsp85_4 sp85_4 sp4_p3 11.551961
Rsn85_4 sn85_4 sn4_p3 11.551961
Rsp85_5 sp85_5 sp5_p3 11.551961
Rsn85_5 sn85_5 sn5_p3 11.551961
Rsp85_6 sp85_6 sp6_p3 11.551961
Rsn85_6 sn85_6 sn6_p3 11.551961
Rsp85_7 sp85_7 sp7_p3 11.551961
Rsn85_7 sn85_7 sn7_p3 11.551961
Rsp85_8 sp85_8 sp8_p3 11.551961
Rsn85_8 sn85_8 sn8_p3 11.551961
Rsp85_9 sp85_9 sp9_p3 11.551961
Rsn85_9 sn85_9 sn9_p3 11.551961
Rsp85_10 sp85_10 sp10_p3 11.551961
Rsn85_10 sn85_10 sn10_p3 11.551961


**********Weight Differntial Op-AMPS and Connecting Resistors****************

XDIFFw1_p1 sp1_p1 sn1_p1 nin1_1 diff3
Rconn1_p1 nin1_1 nin1 1m
XDIFFw2_p1 sp2_p1 sn2_p1 nin2_1 diff3
Rconn2_p1 nin2_1 nin2 1m
XDIFFw3_p1 sp3_p1 sn3_p1 nin3_1 diff3
Rconn3_p1 nin3_1 nin3 1m
XDIFFw4_p1 sp4_p1 sn4_p1 nin4_1 diff3
Rconn4_p1 nin4_1 nin4 1m
XDIFFw5_p1 sp5_p1 sn5_p1 nin5_1 diff3
Rconn5_p1 nin5_1 nin5 1m
XDIFFw6_p1 sp6_p1 sn6_p1 nin6_1 diff3
Rconn6_p1 nin6_1 nin6 1m
XDIFFw7_p1 sp7_p1 sn7_p1 nin7_1 diff3
Rconn7_p1 nin7_1 nin7 1m
XDIFFw8_p1 sp8_p1 sn8_p1 nin8_1 diff3
Rconn8_p1 nin8_1 nin8 1m
XDIFFw9_p1 sp9_p1 sn9_p1 nin9_1 diff3
Rconn9_p1 nin9_1 nin9 1m
XDIFFw10_p1 sp10_p1 sn10_p1 nin10_1 diff3
Rconn10_p1 nin10_1 nin10 1m
XDIFFw1_p2 sp1_p2 sn1_p2 nin1_2 diff3
Rconn1_p2 nin1_2 nin1 1m
XDIFFw2_p2 sp2_p2 sn2_p2 nin2_2 diff3
Rconn2_p2 nin2_2 nin2 1m
XDIFFw3_p2 sp3_p2 sn3_p2 nin3_2 diff3
Rconn3_p2 nin3_2 nin3 1m
XDIFFw4_p2 sp4_p2 sn4_p2 nin4_2 diff3
Rconn4_p2 nin4_2 nin4 1m
XDIFFw5_p2 sp5_p2 sn5_p2 nin5_2 diff3
Rconn5_p2 nin5_2 nin5 1m
XDIFFw6_p2 sp6_p2 sn6_p2 nin6_2 diff3
Rconn6_p2 nin6_2 nin6 1m
XDIFFw7_p2 sp7_p2 sn7_p2 nin7_2 diff3
Rconn7_p2 nin7_2 nin7 1m
XDIFFw8_p2 sp8_p2 sn8_p2 nin8_2 diff3
Rconn8_p2 nin8_2 nin8 1m
XDIFFw9_p2 sp9_p2 sn9_p2 nin9_2 diff3
Rconn9_p2 nin9_2 nin9 1m
XDIFFw10_p2 sp10_p2 sn10_p2 nin10_2 diff3
Rconn10_p2 nin10_2 nin10 1m
XDIFFw1_p3 sp1_p3 sn1_p3 nin1_3 diff3
Rconn1_p3 nin1_3 nin1 1m
XDIFFw2_p3 sp2_p3 sn2_p3 nin2_3 diff3
Rconn2_p3 nin2_3 nin2 1m
XDIFFw3_p3 sp3_p3 sn3_p3 nin3_3 diff3
Rconn3_p3 nin3_3 nin3 1m
XDIFFw4_p3 sp4_p3 sn4_p3 nin4_3 diff3
Rconn4_p3 nin4_3 nin4 1m
XDIFFw5_p3 sp5_p3 sn5_p3 nin5_3 diff3
Rconn5_p3 nin5_3 nin5 1m
XDIFFw6_p3 sp6_p3 sn6_p3 nin6_3 diff3
Rconn6_p3 nin6_3 nin6 1m
XDIFFw7_p3 sp7_p3 sn7_p3 nin7_3 diff3
Rconn7_p3 nin7_3 nin7 1m
XDIFFw8_p3 sp8_p3 sn8_p3 nin8_3 diff3
Rconn8_p3 nin8_3 nin8 1m
XDIFFw9_p3 sp9_p3 sn9_p3 nin9_3 diff3
Rconn9_p3 nin9_3 nin9 1m
XDIFFw10_p3 sp10_p3 sn10_p3 nin10_3 diff3
Rconn10_p3 nin10_3 nin10 1m


**********neurons****************

Xsig1 nin1 out1 vdd 0 neuron
Xsig2 nin2 out2 vdd 0 neuron
Xsig3 nin3 out3 vdd 0 neuron
Xsig4 nin4 out4 vdd 0 neuron
Xsig5 nin5 out5 vdd 0 neuron
Xsig6 nin6 out6 vdd 0 neuron
Xsig7 nin7 out7 vdd 0 neuron
Xsig8 nin8 out8 vdd 0 neuron
Xsig9 nin9 out9 vdd 0 neuron
Xsig10 nin10 out10 vdd 0 neuron
.ENDS layer3