.SUBCKT layer2 vdd vss 0 in1 in2 in3 in4 in5 in6 in7 in8 in9 in10 in11 in12 in13 in14 in15 in16 in17 in18 in19 in20 in21 in22 in23 in24 in25 in26 in27 in28 in29 in30 in31 in32 in33 in34 in35 in36 in37 in38 in39 in40 in41 in42 in43 in44 in45 in46 in47 in48 in49 in50 in51 in52 in53 in54 in55 in56 in57 in58 in59 in60 in61 in62 in63 in64 in65 in66 in67 in68 in69 in70 in71 in72 in73 in74 in75 in76 in77 in78 in79 in80 in81 in82 in83 in84 in85 in86 in87 in88 in89 in90 in91 in92 in93 in94 in95 in96 in97 in98 in99 in100 in101 in102 in103 in104 in105 in106 in107 in108 in109 in110 in111 in112 in113 in114 in115 in116 in117 in118 in119 in120 out1 out2 out3 out4 out5 out6 out7 out8 out9 out10 out11 out12 out13 out14 out15 out16 out17 out18 out19 out20 out21 out22 out23 out24 out25 out26 out27 out28 out29 out30 out31 out32 out33 out34 out35 out36 out37 out38 out39 out40 out41 out42 out43 out44 out45 out46 out47 out48 out49 out50 out51 out52 out53 out54 out55 out56 out57 out58 out59 out60 out61 out62 out63 out64 out65 out66 out67 out68 out69 out70 out71 out72 out73 out74 out75 out76 out77 out78 out79 out80 out81 out82 out83 out84 

**********Positive Weighted Array**********
Rwpos1_1 in1_1 sp1_1 78000.000000
Rwpos1_2 in1_2 sp1_2 202000.000000
Rwpos1_3 in1_3 sp1_3 78000.000000
Rwpos1_4 in1_4 sp1_4 202000.000000
Rwpos1_5 in1_5 sp1_5 202000.000000
Rwpos1_6 in1_6 sp1_6 78000.000000
Rwpos1_7 in1_7 sp1_7 78000.000000
Rwpos1_8 in1_8 sp1_8 202000.000000
Rwpos1_9 in1_9 sp1_9 202000.000000
Rwpos1_10 in1_10 sp1_10 78000.000000
Rwpos1_11 in1_11 sp1_11 78000.000000
Rwpos1_12 in1_12 sp1_12 78000.000000
Rwpos1_13 in1_13 sp1_13 202000.000000
Rwpos1_14 in1_14 sp1_14 202000.000000
Rwpos1_15 in1_15 sp1_15 202000.000000
Rwpos1_16 in1_16 sp1_16 202000.000000
Rwpos1_17 in1_17 sp1_17 78000.000000
Rwpos1_18 in1_18 sp1_18 78000.000000
Rwpos1_19 in1_19 sp1_19 202000.000000
Rwpos1_20 in1_20 sp1_20 202000.000000
Rwpos1_21 in1_21 sp1_21 78000.000000
Rwpos1_22 in1_22 sp1_22 202000.000000
Rwpos1_23 in1_23 sp1_23 78000.000000
Rwpos1_24 in1_24 sp1_24 78000.000000
Rwpos1_25 in1_25 sp1_25 78000.000000
Rwpos1_26 in1_26 sp1_26 78000.000000
Rwpos1_27 in1_27 sp1_27 202000.000000
Rwpos1_28 in1_28 sp1_28 202000.000000
Rwpos1_29 in1_29 sp1_29 202000.000000
Rwpos1_30 in1_30 sp1_30 202000.000000
Rwpos1_31 in1_31 sp1_31 78000.000000
Rwpos1_32 in1_32 sp1_32 78000.000000
Rwpos1_33 in1_33 sp1_33 202000.000000
Rwpos1_34 in1_34 sp1_34 202000.000000
Rwpos1_35 in1_35 sp1_35 78000.000000
Rwpos1_36 in1_36 sp1_36 202000.000000
Rwpos1_37 in1_37 sp1_37 202000.000000
Rwpos1_38 in1_38 sp1_38 202000.000000
Rwpos1_39 in1_39 sp1_39 202000.000000
Rwpos1_40 in1_40 sp1_40 202000.000000
Rwpos1_41 in1_41 sp1_41 202000.000000
Rwpos1_42 in1_42 sp1_42 78000.000000
Rwpos1_43 in1_43 sp1_43 78000.000000
Rwpos1_44 in1_44 sp1_44 202000.000000
Rwpos1_45 in1_45 sp1_45 202000.000000
Rwpos1_46 in1_46 sp1_46 202000.000000
Rwpos1_47 in1_47 sp1_47 78000.000000
Rwpos1_48 in1_48 sp1_48 202000.000000
Rwpos1_49 in1_49 sp1_49 202000.000000
Rwpos1_50 in1_50 sp1_50 202000.000000
Rwpos1_51 in1_51 sp1_51 78000.000000
Rwpos1_52 in1_52 sp1_52 202000.000000
Rwpos1_53 in1_53 sp1_53 202000.000000
Rwpos1_54 in1_54 sp1_54 78000.000000
Rwpos1_55 in1_55 sp1_55 78000.000000
Rwpos1_56 in1_56 sp1_56 78000.000000
Rwpos1_57 in1_57 sp1_57 78000.000000
Rwpos1_58 in1_58 sp1_58 202000.000000
Rwpos1_59 in1_59 sp1_59 78000.000000
Rwpos1_60 in1_60 sp1_60 78000.000000
Rwpos1_61 in1_61 sp1_61 202000.000000
Rwpos1_62 in1_62 sp1_62 78000.000000
Rwpos1_63 in1_63 sp1_63 78000.000000
Rwpos1_64 in1_64 sp1_64 78000.000000
Rwpos1_65 in1_65 sp1_65 78000.000000
Rwpos1_66 in1_66 sp1_66 78000.000000
Rwpos1_67 in1_67 sp1_67 202000.000000
Rwpos1_68 in1_68 sp1_68 78000.000000
Rwpos1_69 in1_69 sp1_69 78000.000000
Rwpos1_70 in1_70 sp1_70 202000.000000
Rwpos1_71 in1_71 sp1_71 78000.000000
Rwpos1_72 in1_72 sp1_72 202000.000000
Rwpos1_73 in1_73 sp1_73 78000.000000
Rwpos1_74 in1_74 sp1_74 202000.000000
Rwpos1_75 in1_75 sp1_75 78000.000000
Rwpos1_76 in1_76 sp1_76 202000.000000
Rwpos1_77 in1_77 sp1_77 78000.000000
Rwpos1_78 in1_78 sp1_78 78000.000000
Rwpos1_79 in1_79 sp1_79 78000.000000
Rwpos1_80 in1_80 sp1_80 78000.000000
Rwpos1_81 in1_81 sp1_81 78000.000000
Rwpos1_82 in1_82 sp1_82 202000.000000
Rwpos1_83 in1_83 sp1_83 78000.000000
Rwpos1_84 in1_84 sp1_84 78000.000000
Rwpos2_1 in2_1 sp2_1 78000.000000
Rwpos2_2 in2_2 sp2_2 78000.000000
Rwpos2_3 in2_3 sp2_3 202000.000000
Rwpos2_4 in2_4 sp2_4 78000.000000
Rwpos2_5 in2_5 sp2_5 78000.000000
Rwpos2_6 in2_6 sp2_6 78000.000000
Rwpos2_7 in2_7 sp2_7 202000.000000
Rwpos2_8 in2_8 sp2_8 78000.000000
Rwpos2_9 in2_9 sp2_9 202000.000000
Rwpos2_10 in2_10 sp2_10 78000.000000
Rwpos2_11 in2_11 sp2_11 78000.000000
Rwpos2_12 in2_12 sp2_12 202000.000000
Rwpos2_13 in2_13 sp2_13 78000.000000
Rwpos2_14 in2_14 sp2_14 78000.000000
Rwpos2_15 in2_15 sp2_15 202000.000000
Rwpos2_16 in2_16 sp2_16 202000.000000
Rwpos2_17 in2_17 sp2_17 78000.000000
Rwpos2_18 in2_18 sp2_18 78000.000000
Rwpos2_19 in2_19 sp2_19 202000.000000
Rwpos2_20 in2_20 sp2_20 202000.000000
Rwpos2_21 in2_21 sp2_21 78000.000000
Rwpos2_22 in2_22 sp2_22 78000.000000
Rwpos2_23 in2_23 sp2_23 78000.000000
Rwpos2_24 in2_24 sp2_24 78000.000000
Rwpos2_25 in2_25 sp2_25 202000.000000
Rwpos2_26 in2_26 sp2_26 78000.000000
Rwpos2_27 in2_27 sp2_27 202000.000000
Rwpos2_28 in2_28 sp2_28 202000.000000
Rwpos2_29 in2_29 sp2_29 78000.000000
Rwpos2_30 in2_30 sp2_30 78000.000000
Rwpos2_31 in2_31 sp2_31 202000.000000
Rwpos2_32 in2_32 sp2_32 202000.000000
Rwpos2_33 in2_33 sp2_33 202000.000000
Rwpos2_34 in2_34 sp2_34 202000.000000
Rwpos2_35 in2_35 sp2_35 202000.000000
Rwpos2_36 in2_36 sp2_36 202000.000000
Rwpos2_37 in2_37 sp2_37 202000.000000
Rwpos2_38 in2_38 sp2_38 202000.000000
Rwpos2_39 in2_39 sp2_39 78000.000000
Rwpos2_40 in2_40 sp2_40 202000.000000
Rwpos2_41 in2_41 sp2_41 202000.000000
Rwpos2_42 in2_42 sp2_42 202000.000000
Rwpos2_43 in2_43 sp2_43 78000.000000
Rwpos2_44 in2_44 sp2_44 78000.000000
Rwpos2_45 in2_45 sp2_45 78000.000000
Rwpos2_46 in2_46 sp2_46 202000.000000
Rwpos2_47 in2_47 sp2_47 78000.000000
Rwpos2_48 in2_48 sp2_48 202000.000000
Rwpos2_49 in2_49 sp2_49 202000.000000
Rwpos2_50 in2_50 sp2_50 202000.000000
Rwpos2_51 in2_51 sp2_51 202000.000000
Rwpos2_52 in2_52 sp2_52 202000.000000
Rwpos2_53 in2_53 sp2_53 78000.000000
Rwpos2_54 in2_54 sp2_54 202000.000000
Rwpos2_55 in2_55 sp2_55 78000.000000
Rwpos2_56 in2_56 sp2_56 78000.000000
Rwpos2_57 in2_57 sp2_57 78000.000000
Rwpos2_58 in2_58 sp2_58 78000.000000
Rwpos2_59 in2_59 sp2_59 202000.000000
Rwpos2_60 in2_60 sp2_60 78000.000000
Rwpos2_61 in2_61 sp2_61 78000.000000
Rwpos2_62 in2_62 sp2_62 78000.000000
Rwpos2_63 in2_63 sp2_63 78000.000000
Rwpos2_64 in2_64 sp2_64 202000.000000
Rwpos2_65 in2_65 sp2_65 78000.000000
Rwpos2_66 in2_66 sp2_66 202000.000000
Rwpos2_67 in2_67 sp2_67 202000.000000
Rwpos2_68 in2_68 sp2_68 78000.000000
Rwpos2_69 in2_69 sp2_69 78000.000000
Rwpos2_70 in2_70 sp2_70 78000.000000
Rwpos2_71 in2_71 sp2_71 78000.000000
Rwpos2_72 in2_72 sp2_72 78000.000000
Rwpos2_73 in2_73 sp2_73 78000.000000
Rwpos2_74 in2_74 sp2_74 78000.000000
Rwpos2_75 in2_75 sp2_75 202000.000000
Rwpos2_76 in2_76 sp2_76 202000.000000
Rwpos2_77 in2_77 sp2_77 202000.000000
Rwpos2_78 in2_78 sp2_78 202000.000000
Rwpos2_79 in2_79 sp2_79 78000.000000
Rwpos2_80 in2_80 sp2_80 78000.000000
Rwpos2_81 in2_81 sp2_81 78000.000000
Rwpos2_82 in2_82 sp2_82 78000.000000
Rwpos2_83 in2_83 sp2_83 78000.000000
Rwpos2_84 in2_84 sp2_84 78000.000000
Rwpos3_1 in3_1 sp3_1 202000.000000
Rwpos3_2 in3_2 sp3_2 202000.000000
Rwpos3_3 in3_3 sp3_3 202000.000000
Rwpos3_4 in3_4 sp3_4 78000.000000
Rwpos3_5 in3_5 sp3_5 202000.000000
Rwpos3_6 in3_6 sp3_6 78000.000000
Rwpos3_7 in3_7 sp3_7 78000.000000
Rwpos3_8 in3_8 sp3_8 202000.000000
Rwpos3_9 in3_9 sp3_9 202000.000000
Rwpos3_10 in3_10 sp3_10 78000.000000
Rwpos3_11 in3_11 sp3_11 78000.000000
Rwpos3_12 in3_12 sp3_12 78000.000000
Rwpos3_13 in3_13 sp3_13 78000.000000
Rwpos3_14 in3_14 sp3_14 78000.000000
Rwpos3_15 in3_15 sp3_15 78000.000000
Rwpos3_16 in3_16 sp3_16 78000.000000
Rwpos3_17 in3_17 sp3_17 202000.000000
Rwpos3_18 in3_18 sp3_18 78000.000000
Rwpos3_19 in3_19 sp3_19 78000.000000
Rwpos3_20 in3_20 sp3_20 78000.000000
Rwpos3_21 in3_21 sp3_21 202000.000000
Rwpos3_22 in3_22 sp3_22 202000.000000
Rwpos3_23 in3_23 sp3_23 202000.000000
Rwpos3_24 in3_24 sp3_24 78000.000000
Rwpos3_25 in3_25 sp3_25 202000.000000
Rwpos3_26 in3_26 sp3_26 78000.000000
Rwpos3_27 in3_27 sp3_27 78000.000000
Rwpos3_28 in3_28 sp3_28 78000.000000
Rwpos3_29 in3_29 sp3_29 202000.000000
Rwpos3_30 in3_30 sp3_30 202000.000000
Rwpos3_31 in3_31 sp3_31 202000.000000
Rwpos3_32 in3_32 sp3_32 78000.000000
Rwpos3_33 in3_33 sp3_33 202000.000000
Rwpos3_34 in3_34 sp3_34 78000.000000
Rwpos3_35 in3_35 sp3_35 202000.000000
Rwpos3_36 in3_36 sp3_36 78000.000000
Rwpos3_37 in3_37 sp3_37 78000.000000
Rwpos3_38 in3_38 sp3_38 78000.000000
Rwpos3_39 in3_39 sp3_39 78000.000000
Rwpos3_40 in3_40 sp3_40 78000.000000
Rwpos3_41 in3_41 sp3_41 202000.000000
Rwpos3_42 in3_42 sp3_42 202000.000000
Rwpos3_43 in3_43 sp3_43 78000.000000
Rwpos3_44 in3_44 sp3_44 202000.000000
Rwpos3_45 in3_45 sp3_45 78000.000000
Rwpos3_46 in3_46 sp3_46 78000.000000
Rwpos3_47 in3_47 sp3_47 78000.000000
Rwpos3_48 in3_48 sp3_48 202000.000000
Rwpos3_49 in3_49 sp3_49 78000.000000
Rwpos3_50 in3_50 sp3_50 78000.000000
Rwpos3_51 in3_51 sp3_51 78000.000000
Rwpos3_52 in3_52 sp3_52 78000.000000
Rwpos3_53 in3_53 sp3_53 202000.000000
Rwpos3_54 in3_54 sp3_54 78000.000000
Rwpos3_55 in3_55 sp3_55 202000.000000
Rwpos3_56 in3_56 sp3_56 78000.000000
Rwpos3_57 in3_57 sp3_57 78000.000000
Rwpos3_58 in3_58 sp3_58 202000.000000
Rwpos3_59 in3_59 sp3_59 78000.000000
Rwpos3_60 in3_60 sp3_60 78000.000000
Rwpos3_61 in3_61 sp3_61 202000.000000
Rwpos3_62 in3_62 sp3_62 202000.000000
Rwpos3_63 in3_63 sp3_63 78000.000000
Rwpos3_64 in3_64 sp3_64 202000.000000
Rwpos3_65 in3_65 sp3_65 202000.000000
Rwpos3_66 in3_66 sp3_66 202000.000000
Rwpos3_67 in3_67 sp3_67 78000.000000
Rwpos3_68 in3_68 sp3_68 78000.000000
Rwpos3_69 in3_69 sp3_69 78000.000000
Rwpos3_70 in3_70 sp3_70 202000.000000
Rwpos3_71 in3_71 sp3_71 202000.000000
Rwpos3_72 in3_72 sp3_72 78000.000000
Rwpos3_73 in3_73 sp3_73 202000.000000
Rwpos3_74 in3_74 sp3_74 202000.000000
Rwpos3_75 in3_75 sp3_75 78000.000000
Rwpos3_76 in3_76 sp3_76 78000.000000
Rwpos3_77 in3_77 sp3_77 78000.000000
Rwpos3_78 in3_78 sp3_78 78000.000000
Rwpos3_79 in3_79 sp3_79 78000.000000
Rwpos3_80 in3_80 sp3_80 202000.000000
Rwpos3_81 in3_81 sp3_81 202000.000000
Rwpos3_82 in3_82 sp3_82 78000.000000
Rwpos3_83 in3_83 sp3_83 202000.000000
Rwpos3_84 in3_84 sp3_84 202000.000000
Rwpos4_1 in4_1 sp4_1 202000.000000
Rwpos4_2 in4_2 sp4_2 202000.000000
Rwpos4_3 in4_3 sp4_3 202000.000000
Rwpos4_4 in4_4 sp4_4 78000.000000
Rwpos4_5 in4_5 sp4_5 78000.000000
Rwpos4_6 in4_6 sp4_6 78000.000000
Rwpos4_7 in4_7 sp4_7 78000.000000
Rwpos4_8 in4_8 sp4_8 202000.000000
Rwpos4_9 in4_9 sp4_9 78000.000000
Rwpos4_10 in4_10 sp4_10 202000.000000
Rwpos4_11 in4_11 sp4_11 78000.000000
Rwpos4_12 in4_12 sp4_12 202000.000000
Rwpos4_13 in4_13 sp4_13 78000.000000
Rwpos4_14 in4_14 sp4_14 78000.000000
Rwpos4_15 in4_15 sp4_15 78000.000000
Rwpos4_16 in4_16 sp4_16 202000.000000
Rwpos4_17 in4_17 sp4_17 78000.000000
Rwpos4_18 in4_18 sp4_18 78000.000000
Rwpos4_19 in4_19 sp4_19 202000.000000
Rwpos4_20 in4_20 sp4_20 202000.000000
Rwpos4_21 in4_21 sp4_21 78000.000000
Rwpos4_22 in4_22 sp4_22 202000.000000
Rwpos4_23 in4_23 sp4_23 78000.000000
Rwpos4_24 in4_24 sp4_24 78000.000000
Rwpos4_25 in4_25 sp4_25 78000.000000
Rwpos4_26 in4_26 sp4_26 78000.000000
Rwpos4_27 in4_27 sp4_27 78000.000000
Rwpos4_28 in4_28 sp4_28 78000.000000
Rwpos4_29 in4_29 sp4_29 202000.000000
Rwpos4_30 in4_30 sp4_30 78000.000000
Rwpos4_31 in4_31 sp4_31 78000.000000
Rwpos4_32 in4_32 sp4_32 78000.000000
Rwpos4_33 in4_33 sp4_33 202000.000000
Rwpos4_34 in4_34 sp4_34 78000.000000
Rwpos4_35 in4_35 sp4_35 78000.000000
Rwpos4_36 in4_36 sp4_36 202000.000000
Rwpos4_37 in4_37 sp4_37 78000.000000
Rwpos4_38 in4_38 sp4_38 202000.000000
Rwpos4_39 in4_39 sp4_39 78000.000000
Rwpos4_40 in4_40 sp4_40 202000.000000
Rwpos4_41 in4_41 sp4_41 202000.000000
Rwpos4_42 in4_42 sp4_42 78000.000000
Rwpos4_43 in4_43 sp4_43 78000.000000
Rwpos4_44 in4_44 sp4_44 202000.000000
Rwpos4_45 in4_45 sp4_45 202000.000000
Rwpos4_46 in4_46 sp4_46 78000.000000
Rwpos4_47 in4_47 sp4_47 78000.000000
Rwpos4_48 in4_48 sp4_48 202000.000000
Rwpos4_49 in4_49 sp4_49 202000.000000
Rwpos4_50 in4_50 sp4_50 78000.000000
Rwpos4_51 in4_51 sp4_51 78000.000000
Rwpos4_52 in4_52 sp4_52 78000.000000
Rwpos4_53 in4_53 sp4_53 202000.000000
Rwpos4_54 in4_54 sp4_54 78000.000000
Rwpos4_55 in4_55 sp4_55 202000.000000
Rwpos4_56 in4_56 sp4_56 202000.000000
Rwpos4_57 in4_57 sp4_57 202000.000000
Rwpos4_58 in4_58 sp4_58 202000.000000
Rwpos4_59 in4_59 sp4_59 202000.000000
Rwpos4_60 in4_60 sp4_60 78000.000000
Rwpos4_61 in4_61 sp4_61 202000.000000
Rwpos4_62 in4_62 sp4_62 78000.000000
Rwpos4_63 in4_63 sp4_63 202000.000000
Rwpos4_64 in4_64 sp4_64 202000.000000
Rwpos4_65 in4_65 sp4_65 202000.000000
Rwpos4_66 in4_66 sp4_66 202000.000000
Rwpos4_67 in4_67 sp4_67 202000.000000
Rwpos4_68 in4_68 sp4_68 202000.000000
Rwpos4_69 in4_69 sp4_69 202000.000000
Rwpos4_70 in4_70 sp4_70 202000.000000
Rwpos4_71 in4_71 sp4_71 202000.000000
Rwpos4_72 in4_72 sp4_72 202000.000000
Rwpos4_73 in4_73 sp4_73 202000.000000
Rwpos4_74 in4_74 sp4_74 202000.000000
Rwpos4_75 in4_75 sp4_75 202000.000000
Rwpos4_76 in4_76 sp4_76 202000.000000
Rwpos4_77 in4_77 sp4_77 78000.000000
Rwpos4_78 in4_78 sp4_78 78000.000000
Rwpos4_79 in4_79 sp4_79 202000.000000
Rwpos4_80 in4_80 sp4_80 78000.000000
Rwpos4_81 in4_81 sp4_81 78000.000000
Rwpos4_82 in4_82 sp4_82 202000.000000
Rwpos4_83 in4_83 sp4_83 202000.000000
Rwpos4_84 in4_84 sp4_84 202000.000000
Rwpos5_1 in5_1 sp5_1 78000.000000
Rwpos5_2 in5_2 sp5_2 78000.000000
Rwpos5_3 in5_3 sp5_3 202000.000000
Rwpos5_4 in5_4 sp5_4 78000.000000
Rwpos5_5 in5_5 sp5_5 78000.000000
Rwpos5_6 in5_6 sp5_6 78000.000000
Rwpos5_7 in5_7 sp5_7 202000.000000
Rwpos5_8 in5_8 sp5_8 78000.000000
Rwpos5_9 in5_9 sp5_9 78000.000000
Rwpos5_10 in5_10 sp5_10 78000.000000
Rwpos5_11 in5_11 sp5_11 78000.000000
Rwpos5_12 in5_12 sp5_12 78000.000000
Rwpos5_13 in5_13 sp5_13 78000.000000
Rwpos5_14 in5_14 sp5_14 202000.000000
Rwpos5_15 in5_15 sp5_15 78000.000000
Rwpos5_16 in5_16 sp5_16 78000.000000
Rwpos5_17 in5_17 sp5_17 202000.000000
Rwpos5_18 in5_18 sp5_18 78000.000000
Rwpos5_19 in5_19 sp5_19 78000.000000
Rwpos5_20 in5_20 sp5_20 202000.000000
Rwpos5_21 in5_21 sp5_21 202000.000000
Rwpos5_22 in5_22 sp5_22 202000.000000
Rwpos5_23 in5_23 sp5_23 202000.000000
Rwpos5_24 in5_24 sp5_24 78000.000000
Rwpos5_25 in5_25 sp5_25 202000.000000
Rwpos5_26 in5_26 sp5_26 78000.000000
Rwpos5_27 in5_27 sp5_27 78000.000000
Rwpos5_28 in5_28 sp5_28 78000.000000
Rwpos5_29 in5_29 sp5_29 78000.000000
Rwpos5_30 in5_30 sp5_30 78000.000000
Rwpos5_31 in5_31 sp5_31 78000.000000
Rwpos5_32 in5_32 sp5_32 202000.000000
Rwpos5_33 in5_33 sp5_33 202000.000000
Rwpos5_34 in5_34 sp5_34 202000.000000
Rwpos5_35 in5_35 sp5_35 202000.000000
Rwpos5_36 in5_36 sp5_36 202000.000000
Rwpos5_37 in5_37 sp5_37 202000.000000
Rwpos5_38 in5_38 sp5_38 78000.000000
Rwpos5_39 in5_39 sp5_39 202000.000000
Rwpos5_40 in5_40 sp5_40 78000.000000
Rwpos5_41 in5_41 sp5_41 78000.000000
Rwpos5_42 in5_42 sp5_42 78000.000000
Rwpos5_43 in5_43 sp5_43 78000.000000
Rwpos5_44 in5_44 sp5_44 78000.000000
Rwpos5_45 in5_45 sp5_45 202000.000000
Rwpos5_46 in5_46 sp5_46 202000.000000
Rwpos5_47 in5_47 sp5_47 202000.000000
Rwpos5_48 in5_48 sp5_48 202000.000000
Rwpos5_49 in5_49 sp5_49 78000.000000
Rwpos5_50 in5_50 sp5_50 202000.000000
Rwpos5_51 in5_51 sp5_51 78000.000000
Rwpos5_52 in5_52 sp5_52 78000.000000
Rwpos5_53 in5_53 sp5_53 202000.000000
Rwpos5_54 in5_54 sp5_54 78000.000000
Rwpos5_55 in5_55 sp5_55 78000.000000
Rwpos5_56 in5_56 sp5_56 202000.000000
Rwpos5_57 in5_57 sp5_57 202000.000000
Rwpos5_58 in5_58 sp5_58 78000.000000
Rwpos5_59 in5_59 sp5_59 202000.000000
Rwpos5_60 in5_60 sp5_60 78000.000000
Rwpos5_61 in5_61 sp5_61 202000.000000
Rwpos5_62 in5_62 sp5_62 78000.000000
Rwpos5_63 in5_63 sp5_63 202000.000000
Rwpos5_64 in5_64 sp5_64 202000.000000
Rwpos5_65 in5_65 sp5_65 202000.000000
Rwpos5_66 in5_66 sp5_66 78000.000000
Rwpos5_67 in5_67 sp5_67 202000.000000
Rwpos5_68 in5_68 sp5_68 78000.000000
Rwpos5_69 in5_69 sp5_69 202000.000000
Rwpos5_70 in5_70 sp5_70 78000.000000
Rwpos5_71 in5_71 sp5_71 202000.000000
Rwpos5_72 in5_72 sp5_72 202000.000000
Rwpos5_73 in5_73 sp5_73 78000.000000
Rwpos5_74 in5_74 sp5_74 202000.000000
Rwpos5_75 in5_75 sp5_75 202000.000000
Rwpos5_76 in5_76 sp5_76 78000.000000
Rwpos5_77 in5_77 sp5_77 202000.000000
Rwpos5_78 in5_78 sp5_78 78000.000000
Rwpos5_79 in5_79 sp5_79 202000.000000
Rwpos5_80 in5_80 sp5_80 202000.000000
Rwpos5_81 in5_81 sp5_81 202000.000000
Rwpos5_82 in5_82 sp5_82 78000.000000
Rwpos5_83 in5_83 sp5_83 202000.000000
Rwpos5_84 in5_84 sp5_84 78000.000000
Rwpos6_1 in6_1 sp6_1 202000.000000
Rwpos6_2 in6_2 sp6_2 78000.000000
Rwpos6_3 in6_3 sp6_3 202000.000000
Rwpos6_4 in6_4 sp6_4 78000.000000
Rwpos6_5 in6_5 sp6_5 202000.000000
Rwpos6_6 in6_6 sp6_6 78000.000000
Rwpos6_7 in6_7 sp6_7 202000.000000
Rwpos6_8 in6_8 sp6_8 202000.000000
Rwpos6_9 in6_9 sp6_9 78000.000000
Rwpos6_10 in6_10 sp6_10 78000.000000
Rwpos6_11 in6_11 sp6_11 202000.000000
Rwpos6_12 in6_12 sp6_12 78000.000000
Rwpos6_13 in6_13 sp6_13 202000.000000
Rwpos6_14 in6_14 sp6_14 202000.000000
Rwpos6_15 in6_15 sp6_15 202000.000000
Rwpos6_16 in6_16 sp6_16 78000.000000
Rwpos6_17 in6_17 sp6_17 202000.000000
Rwpos6_18 in6_18 sp6_18 202000.000000
Rwpos6_19 in6_19 sp6_19 78000.000000
Rwpos6_20 in6_20 sp6_20 78000.000000
Rwpos6_21 in6_21 sp6_21 202000.000000
Rwpos6_22 in6_22 sp6_22 202000.000000
Rwpos6_23 in6_23 sp6_23 202000.000000
Rwpos6_24 in6_24 sp6_24 202000.000000
Rwpos6_25 in6_25 sp6_25 202000.000000
Rwpos6_26 in6_26 sp6_26 202000.000000
Rwpos6_27 in6_27 sp6_27 202000.000000
Rwpos6_28 in6_28 sp6_28 78000.000000
Rwpos6_29 in6_29 sp6_29 78000.000000
Rwpos6_30 in6_30 sp6_30 78000.000000
Rwpos6_31 in6_31 sp6_31 202000.000000
Rwpos6_32 in6_32 sp6_32 202000.000000
Rwpos6_33 in6_33 sp6_33 78000.000000
Rwpos6_34 in6_34 sp6_34 78000.000000
Rwpos6_35 in6_35 sp6_35 78000.000000
Rwpos6_36 in6_36 sp6_36 202000.000000
Rwpos6_37 in6_37 sp6_37 202000.000000
Rwpos6_38 in6_38 sp6_38 78000.000000
Rwpos6_39 in6_39 sp6_39 202000.000000
Rwpos6_40 in6_40 sp6_40 78000.000000
Rwpos6_41 in6_41 sp6_41 202000.000000
Rwpos6_42 in6_42 sp6_42 202000.000000
Rwpos6_43 in6_43 sp6_43 78000.000000
Rwpos6_44 in6_44 sp6_44 202000.000000
Rwpos6_45 in6_45 sp6_45 78000.000000
Rwpos6_46 in6_46 sp6_46 202000.000000
Rwpos6_47 in6_47 sp6_47 78000.000000
Rwpos6_48 in6_48 sp6_48 202000.000000
Rwpos6_49 in6_49 sp6_49 78000.000000
Rwpos6_50 in6_50 sp6_50 202000.000000
Rwpos6_51 in6_51 sp6_51 202000.000000
Rwpos6_52 in6_52 sp6_52 78000.000000
Rwpos6_53 in6_53 sp6_53 78000.000000
Rwpos6_54 in6_54 sp6_54 202000.000000
Rwpos6_55 in6_55 sp6_55 78000.000000
Rwpos6_56 in6_56 sp6_56 202000.000000
Rwpos6_57 in6_57 sp6_57 202000.000000
Rwpos6_58 in6_58 sp6_58 202000.000000
Rwpos6_59 in6_59 sp6_59 202000.000000
Rwpos6_60 in6_60 sp6_60 78000.000000
Rwpos6_61 in6_61 sp6_61 78000.000000
Rwpos6_62 in6_62 sp6_62 202000.000000
Rwpos6_63 in6_63 sp6_63 78000.000000
Rwpos6_64 in6_64 sp6_64 202000.000000
Rwpos6_65 in6_65 sp6_65 78000.000000
Rwpos6_66 in6_66 sp6_66 202000.000000
Rwpos6_67 in6_67 sp6_67 78000.000000
Rwpos6_68 in6_68 sp6_68 202000.000000
Rwpos6_69 in6_69 sp6_69 202000.000000
Rwpos6_70 in6_70 sp6_70 78000.000000
Rwpos6_71 in6_71 sp6_71 202000.000000
Rwpos6_72 in6_72 sp6_72 78000.000000
Rwpos6_73 in6_73 sp6_73 202000.000000
Rwpos6_74 in6_74 sp6_74 202000.000000
Rwpos6_75 in6_75 sp6_75 78000.000000
Rwpos6_76 in6_76 sp6_76 78000.000000
Rwpos6_77 in6_77 sp6_77 78000.000000
Rwpos6_78 in6_78 sp6_78 78000.000000
Rwpos6_79 in6_79 sp6_79 202000.000000
Rwpos6_80 in6_80 sp6_80 202000.000000
Rwpos6_81 in6_81 sp6_81 202000.000000
Rwpos6_82 in6_82 sp6_82 202000.000000
Rwpos6_83 in6_83 sp6_83 202000.000000
Rwpos6_84 in6_84 sp6_84 202000.000000
Rwpos7_1 in7_1 sp7_1 78000.000000
Rwpos7_2 in7_2 sp7_2 202000.000000
Rwpos7_3 in7_3 sp7_3 202000.000000
Rwpos7_4 in7_4 sp7_4 202000.000000
Rwpos7_5 in7_5 sp7_5 78000.000000
Rwpos7_6 in7_6 sp7_6 78000.000000
Rwpos7_7 in7_7 sp7_7 78000.000000
Rwpos7_8 in7_8 sp7_8 202000.000000
Rwpos7_9 in7_9 sp7_9 78000.000000
Rwpos7_10 in7_10 sp7_10 78000.000000
Rwpos7_11 in7_11 sp7_11 202000.000000
Rwpos7_12 in7_12 sp7_12 78000.000000
Rwpos7_13 in7_13 sp7_13 202000.000000
Rwpos7_14 in7_14 sp7_14 78000.000000
Rwpos7_15 in7_15 sp7_15 202000.000000
Rwpos7_16 in7_16 sp7_16 202000.000000
Rwpos7_17 in7_17 sp7_17 78000.000000
Rwpos7_18 in7_18 sp7_18 78000.000000
Rwpos7_19 in7_19 sp7_19 202000.000000
Rwpos7_20 in7_20 sp7_20 202000.000000
Rwpos7_21 in7_21 sp7_21 202000.000000
Rwpos7_22 in7_22 sp7_22 202000.000000
Rwpos7_23 in7_23 sp7_23 202000.000000
Rwpos7_24 in7_24 sp7_24 78000.000000
Rwpos7_25 in7_25 sp7_25 78000.000000
Rwpos7_26 in7_26 sp7_26 202000.000000
Rwpos7_27 in7_27 sp7_27 78000.000000
Rwpos7_28 in7_28 sp7_28 78000.000000
Rwpos7_29 in7_29 sp7_29 78000.000000
Rwpos7_30 in7_30 sp7_30 78000.000000
Rwpos7_31 in7_31 sp7_31 202000.000000
Rwpos7_32 in7_32 sp7_32 78000.000000
Rwpos7_33 in7_33 sp7_33 202000.000000
Rwpos7_34 in7_34 sp7_34 78000.000000
Rwpos7_35 in7_35 sp7_35 202000.000000
Rwpos7_36 in7_36 sp7_36 78000.000000
Rwpos7_37 in7_37 sp7_37 202000.000000
Rwpos7_38 in7_38 sp7_38 78000.000000
Rwpos7_39 in7_39 sp7_39 78000.000000
Rwpos7_40 in7_40 sp7_40 202000.000000
Rwpos7_41 in7_41 sp7_41 202000.000000
Rwpos7_42 in7_42 sp7_42 78000.000000
Rwpos7_43 in7_43 sp7_43 78000.000000
Rwpos7_44 in7_44 sp7_44 78000.000000
Rwpos7_45 in7_45 sp7_45 202000.000000
Rwpos7_46 in7_46 sp7_46 78000.000000
Rwpos7_47 in7_47 sp7_47 78000.000000
Rwpos7_48 in7_48 sp7_48 202000.000000
Rwpos7_49 in7_49 sp7_49 78000.000000
Rwpos7_50 in7_50 sp7_50 202000.000000
Rwpos7_51 in7_51 sp7_51 202000.000000
Rwpos7_52 in7_52 sp7_52 78000.000000
Rwpos7_53 in7_53 sp7_53 78000.000000
Rwpos7_54 in7_54 sp7_54 202000.000000
Rwpos7_55 in7_55 sp7_55 202000.000000
Rwpos7_56 in7_56 sp7_56 202000.000000
Rwpos7_57 in7_57 sp7_57 202000.000000
Rwpos7_58 in7_58 sp7_58 202000.000000
Rwpos7_59 in7_59 sp7_59 202000.000000
Rwpos7_60 in7_60 sp7_60 78000.000000
Rwpos7_61 in7_61 sp7_61 202000.000000
Rwpos7_62 in7_62 sp7_62 78000.000000
Rwpos7_63 in7_63 sp7_63 78000.000000
Rwpos7_64 in7_64 sp7_64 78000.000000
Rwpos7_65 in7_65 sp7_65 78000.000000
Rwpos7_66 in7_66 sp7_66 78000.000000
Rwpos7_67 in7_67 sp7_67 78000.000000
Rwpos7_68 in7_68 sp7_68 78000.000000
Rwpos7_69 in7_69 sp7_69 78000.000000
Rwpos7_70 in7_70 sp7_70 78000.000000
Rwpos7_71 in7_71 sp7_71 78000.000000
Rwpos7_72 in7_72 sp7_72 78000.000000
Rwpos7_73 in7_73 sp7_73 202000.000000
Rwpos7_74 in7_74 sp7_74 78000.000000
Rwpos7_75 in7_75 sp7_75 202000.000000
Rwpos7_76 in7_76 sp7_76 78000.000000
Rwpos7_77 in7_77 sp7_77 78000.000000
Rwpos7_78 in7_78 sp7_78 78000.000000
Rwpos7_79 in7_79 sp7_79 78000.000000
Rwpos7_80 in7_80 sp7_80 202000.000000
Rwpos7_81 in7_81 sp7_81 202000.000000
Rwpos7_82 in7_82 sp7_82 78000.000000
Rwpos7_83 in7_83 sp7_83 202000.000000
Rwpos7_84 in7_84 sp7_84 202000.000000
Rwpos8_1 in8_1 sp8_1 202000.000000
Rwpos8_2 in8_2 sp8_2 78000.000000
Rwpos8_3 in8_3 sp8_3 78000.000000
Rwpos8_4 in8_4 sp8_4 202000.000000
Rwpos8_5 in8_5 sp8_5 202000.000000
Rwpos8_6 in8_6 sp8_6 78000.000000
Rwpos8_7 in8_7 sp8_7 78000.000000
Rwpos8_8 in8_8 sp8_8 202000.000000
Rwpos8_9 in8_9 sp8_9 202000.000000
Rwpos8_10 in8_10 sp8_10 202000.000000
Rwpos8_11 in8_11 sp8_11 202000.000000
Rwpos8_12 in8_12 sp8_12 202000.000000
Rwpos8_13 in8_13 sp8_13 202000.000000
Rwpos8_14 in8_14 sp8_14 78000.000000
Rwpos8_15 in8_15 sp8_15 202000.000000
Rwpos8_16 in8_16 sp8_16 202000.000000
Rwpos8_17 in8_17 sp8_17 78000.000000
Rwpos8_18 in8_18 sp8_18 202000.000000
Rwpos8_19 in8_19 sp8_19 202000.000000
Rwpos8_20 in8_20 sp8_20 202000.000000
Rwpos8_21 in8_21 sp8_21 202000.000000
Rwpos8_22 in8_22 sp8_22 202000.000000
Rwpos8_23 in8_23 sp8_23 78000.000000
Rwpos8_24 in8_24 sp8_24 78000.000000
Rwpos8_25 in8_25 sp8_25 202000.000000
Rwpos8_26 in8_26 sp8_26 78000.000000
Rwpos8_27 in8_27 sp8_27 202000.000000
Rwpos8_28 in8_28 sp8_28 202000.000000
Rwpos8_29 in8_29 sp8_29 202000.000000
Rwpos8_30 in8_30 sp8_30 78000.000000
Rwpos8_31 in8_31 sp8_31 78000.000000
Rwpos8_32 in8_32 sp8_32 202000.000000
Rwpos8_33 in8_33 sp8_33 78000.000000
Rwpos8_34 in8_34 sp8_34 202000.000000
Rwpos8_35 in8_35 sp8_35 202000.000000
Rwpos8_36 in8_36 sp8_36 202000.000000
Rwpos8_37 in8_37 sp8_37 78000.000000
Rwpos8_38 in8_38 sp8_38 202000.000000
Rwpos8_39 in8_39 sp8_39 202000.000000
Rwpos8_40 in8_40 sp8_40 78000.000000
Rwpos8_41 in8_41 sp8_41 78000.000000
Rwpos8_42 in8_42 sp8_42 78000.000000
Rwpos8_43 in8_43 sp8_43 78000.000000
Rwpos8_44 in8_44 sp8_44 78000.000000
Rwpos8_45 in8_45 sp8_45 202000.000000
Rwpos8_46 in8_46 sp8_46 78000.000000
Rwpos8_47 in8_47 sp8_47 78000.000000
Rwpos8_48 in8_48 sp8_48 202000.000000
Rwpos8_49 in8_49 sp8_49 78000.000000
Rwpos8_50 in8_50 sp8_50 202000.000000
Rwpos8_51 in8_51 sp8_51 78000.000000
Rwpos8_52 in8_52 sp8_52 202000.000000
Rwpos8_53 in8_53 sp8_53 202000.000000
Rwpos8_54 in8_54 sp8_54 202000.000000
Rwpos8_55 in8_55 sp8_55 202000.000000
Rwpos8_56 in8_56 sp8_56 202000.000000
Rwpos8_57 in8_57 sp8_57 78000.000000
Rwpos8_58 in8_58 sp8_58 78000.000000
Rwpos8_59 in8_59 sp8_59 78000.000000
Rwpos8_60 in8_60 sp8_60 78000.000000
Rwpos8_61 in8_61 sp8_61 78000.000000
Rwpos8_62 in8_62 sp8_62 202000.000000
Rwpos8_63 in8_63 sp8_63 202000.000000
Rwpos8_64 in8_64 sp8_64 202000.000000
Rwpos8_65 in8_65 sp8_65 78000.000000
Rwpos8_66 in8_66 sp8_66 202000.000000
Rwpos8_67 in8_67 sp8_67 78000.000000
Rwpos8_68 in8_68 sp8_68 202000.000000
Rwpos8_69 in8_69 sp8_69 78000.000000
Rwpos8_70 in8_70 sp8_70 202000.000000
Rwpos8_71 in8_71 sp8_71 202000.000000
Rwpos8_72 in8_72 sp8_72 78000.000000
Rwpos8_73 in8_73 sp8_73 78000.000000
Rwpos8_74 in8_74 sp8_74 202000.000000
Rwpos8_75 in8_75 sp8_75 78000.000000
Rwpos8_76 in8_76 sp8_76 202000.000000
Rwpos8_77 in8_77 sp8_77 78000.000000
Rwpos8_78 in8_78 sp8_78 202000.000000
Rwpos8_79 in8_79 sp8_79 78000.000000
Rwpos8_80 in8_80 sp8_80 202000.000000
Rwpos8_81 in8_81 sp8_81 78000.000000
Rwpos8_82 in8_82 sp8_82 202000.000000
Rwpos8_83 in8_83 sp8_83 78000.000000
Rwpos8_84 in8_84 sp8_84 202000.000000
Rwpos9_1 in9_1 sp9_1 78000.000000
Rwpos9_2 in9_2 sp9_2 78000.000000
Rwpos9_3 in9_3 sp9_3 78000.000000
Rwpos9_4 in9_4 sp9_4 78000.000000
Rwpos9_5 in9_5 sp9_5 202000.000000
Rwpos9_6 in9_6 sp9_6 78000.000000
Rwpos9_7 in9_7 sp9_7 78000.000000
Rwpos9_8 in9_8 sp9_8 202000.000000
Rwpos9_9 in9_9 sp9_9 78000.000000
Rwpos9_10 in9_10 sp9_10 78000.000000
Rwpos9_11 in9_11 sp9_11 78000.000000
Rwpos9_12 in9_12 sp9_12 78000.000000
Rwpos9_13 in9_13 sp9_13 202000.000000
Rwpos9_14 in9_14 sp9_14 202000.000000
Rwpos9_15 in9_15 sp9_15 78000.000000
Rwpos9_16 in9_16 sp9_16 202000.000000
Rwpos9_17 in9_17 sp9_17 202000.000000
Rwpos9_18 in9_18 sp9_18 202000.000000
Rwpos9_19 in9_19 sp9_19 202000.000000
Rwpos9_20 in9_20 sp9_20 78000.000000
Rwpos9_21 in9_21 sp9_21 78000.000000
Rwpos9_22 in9_22 sp9_22 78000.000000
Rwpos9_23 in9_23 sp9_23 202000.000000
Rwpos9_24 in9_24 sp9_24 78000.000000
Rwpos9_25 in9_25 sp9_25 78000.000000
Rwpos9_26 in9_26 sp9_26 78000.000000
Rwpos9_27 in9_27 sp9_27 202000.000000
Rwpos9_28 in9_28 sp9_28 202000.000000
Rwpos9_29 in9_29 sp9_29 202000.000000
Rwpos9_30 in9_30 sp9_30 78000.000000
Rwpos9_31 in9_31 sp9_31 78000.000000
Rwpos9_32 in9_32 sp9_32 78000.000000
Rwpos9_33 in9_33 sp9_33 78000.000000
Rwpos9_34 in9_34 sp9_34 202000.000000
Rwpos9_35 in9_35 sp9_35 78000.000000
Rwpos9_36 in9_36 sp9_36 78000.000000
Rwpos9_37 in9_37 sp9_37 78000.000000
Rwpos9_38 in9_38 sp9_38 78000.000000
Rwpos9_39 in9_39 sp9_39 202000.000000
Rwpos9_40 in9_40 sp9_40 202000.000000
Rwpos9_41 in9_41 sp9_41 78000.000000
Rwpos9_42 in9_42 sp9_42 78000.000000
Rwpos9_43 in9_43 sp9_43 78000.000000
Rwpos9_44 in9_44 sp9_44 202000.000000
Rwpos9_45 in9_45 sp9_45 78000.000000
Rwpos9_46 in9_46 sp9_46 78000.000000
Rwpos9_47 in9_47 sp9_47 202000.000000
Rwpos9_48 in9_48 sp9_48 78000.000000
Rwpos9_49 in9_49 sp9_49 78000.000000
Rwpos9_50 in9_50 sp9_50 78000.000000
Rwpos9_51 in9_51 sp9_51 202000.000000
Rwpos9_52 in9_52 sp9_52 78000.000000
Rwpos9_53 in9_53 sp9_53 78000.000000
Rwpos9_54 in9_54 sp9_54 202000.000000
Rwpos9_55 in9_55 sp9_55 202000.000000
Rwpos9_56 in9_56 sp9_56 78000.000000
Rwpos9_57 in9_57 sp9_57 78000.000000
Rwpos9_58 in9_58 sp9_58 202000.000000
Rwpos9_59 in9_59 sp9_59 78000.000000
Rwpos9_60 in9_60 sp9_60 78000.000000
Rwpos9_61 in9_61 sp9_61 78000.000000
Rwpos9_62 in9_62 sp9_62 202000.000000
Rwpos9_63 in9_63 sp9_63 78000.000000
Rwpos9_64 in9_64 sp9_64 202000.000000
Rwpos9_65 in9_65 sp9_65 78000.000000
Rwpos9_66 in9_66 sp9_66 78000.000000
Rwpos9_67 in9_67 sp9_67 202000.000000
Rwpos9_68 in9_68 sp9_68 202000.000000
Rwpos9_69 in9_69 sp9_69 202000.000000
Rwpos9_70 in9_70 sp9_70 78000.000000
Rwpos9_71 in9_71 sp9_71 78000.000000
Rwpos9_72 in9_72 sp9_72 78000.000000
Rwpos9_73 in9_73 sp9_73 78000.000000
Rwpos9_74 in9_74 sp9_74 78000.000000
Rwpos9_75 in9_75 sp9_75 78000.000000
Rwpos9_76 in9_76 sp9_76 78000.000000
Rwpos9_77 in9_77 sp9_77 202000.000000
Rwpos9_78 in9_78 sp9_78 78000.000000
Rwpos9_79 in9_79 sp9_79 78000.000000
Rwpos9_80 in9_80 sp9_80 202000.000000
Rwpos9_81 in9_81 sp9_81 202000.000000
Rwpos9_82 in9_82 sp9_82 78000.000000
Rwpos9_83 in9_83 sp9_83 202000.000000
Rwpos9_84 in9_84 sp9_84 78000.000000
Rwpos10_1 in10_1 sp10_1 78000.000000
Rwpos10_2 in10_2 sp10_2 202000.000000
Rwpos10_3 in10_3 sp10_3 202000.000000
Rwpos10_4 in10_4 sp10_4 78000.000000
Rwpos10_5 in10_5 sp10_5 202000.000000
Rwpos10_6 in10_6 sp10_6 78000.000000
Rwpos10_7 in10_7 sp10_7 78000.000000
Rwpos10_8 in10_8 sp10_8 202000.000000
Rwpos10_9 in10_9 sp10_9 78000.000000
Rwpos10_10 in10_10 sp10_10 202000.000000
Rwpos10_11 in10_11 sp10_11 78000.000000
Rwpos10_12 in10_12 sp10_12 202000.000000
Rwpos10_13 in10_13 sp10_13 78000.000000
Rwpos10_14 in10_14 sp10_14 78000.000000
Rwpos10_15 in10_15 sp10_15 202000.000000
Rwpos10_16 in10_16 sp10_16 78000.000000
Rwpos10_17 in10_17 sp10_17 78000.000000
Rwpos10_18 in10_18 sp10_18 202000.000000
Rwpos10_19 in10_19 sp10_19 78000.000000
Rwpos10_20 in10_20 sp10_20 78000.000000
Rwpos10_21 in10_21 sp10_21 202000.000000
Rwpos10_22 in10_22 sp10_22 202000.000000
Rwpos10_23 in10_23 sp10_23 202000.000000
Rwpos10_24 in10_24 sp10_24 202000.000000
Rwpos10_25 in10_25 sp10_25 78000.000000
Rwpos10_26 in10_26 sp10_26 202000.000000
Rwpos10_27 in10_27 sp10_27 78000.000000
Rwpos10_28 in10_28 sp10_28 78000.000000
Rwpos10_29 in10_29 sp10_29 202000.000000
Rwpos10_30 in10_30 sp10_30 78000.000000
Rwpos10_31 in10_31 sp10_31 78000.000000
Rwpos10_32 in10_32 sp10_32 202000.000000
Rwpos10_33 in10_33 sp10_33 202000.000000
Rwpos10_34 in10_34 sp10_34 78000.000000
Rwpos10_35 in10_35 sp10_35 202000.000000
Rwpos10_36 in10_36 sp10_36 202000.000000
Rwpos10_37 in10_37 sp10_37 78000.000000
Rwpos10_38 in10_38 sp10_38 78000.000000
Rwpos10_39 in10_39 sp10_39 78000.000000
Rwpos10_40 in10_40 sp10_40 78000.000000
Rwpos10_41 in10_41 sp10_41 202000.000000
Rwpos10_42 in10_42 sp10_42 202000.000000
Rwpos10_43 in10_43 sp10_43 78000.000000
Rwpos10_44 in10_44 sp10_44 202000.000000
Rwpos10_45 in10_45 sp10_45 202000.000000
Rwpos10_46 in10_46 sp10_46 78000.000000
Rwpos10_47 in10_47 sp10_47 78000.000000
Rwpos10_48 in10_48 sp10_48 78000.000000
Rwpos10_49 in10_49 sp10_49 78000.000000
Rwpos10_50 in10_50 sp10_50 78000.000000
Rwpos10_51 in10_51 sp10_51 78000.000000
Rwpos10_52 in10_52 sp10_52 78000.000000
Rwpos10_53 in10_53 sp10_53 78000.000000
Rwpos10_54 in10_54 sp10_54 78000.000000
Rwpos10_55 in10_55 sp10_55 78000.000000
Rwpos10_56 in10_56 sp10_56 202000.000000
Rwpos10_57 in10_57 sp10_57 202000.000000
Rwpos10_58 in10_58 sp10_58 202000.000000
Rwpos10_59 in10_59 sp10_59 202000.000000
Rwpos10_60 in10_60 sp10_60 202000.000000
Rwpos10_61 in10_61 sp10_61 202000.000000
Rwpos10_62 in10_62 sp10_62 78000.000000
Rwpos10_63 in10_63 sp10_63 202000.000000
Rwpos10_64 in10_64 sp10_64 78000.000000
Rwpos10_65 in10_65 sp10_65 202000.000000
Rwpos10_66 in10_66 sp10_66 202000.000000
Rwpos10_67 in10_67 sp10_67 78000.000000
Rwpos10_68 in10_68 sp10_68 78000.000000
Rwpos10_69 in10_69 sp10_69 202000.000000
Rwpos10_70 in10_70 sp10_70 202000.000000
Rwpos10_71 in10_71 sp10_71 202000.000000
Rwpos10_72 in10_72 sp10_72 202000.000000
Rwpos10_73 in10_73 sp10_73 202000.000000
Rwpos10_74 in10_74 sp10_74 78000.000000
Rwpos10_75 in10_75 sp10_75 202000.000000
Rwpos10_76 in10_76 sp10_76 202000.000000
Rwpos10_77 in10_77 sp10_77 202000.000000
Rwpos10_78 in10_78 sp10_78 202000.000000
Rwpos10_79 in10_79 sp10_79 78000.000000
Rwpos10_80 in10_80 sp10_80 202000.000000
Rwpos10_81 in10_81 sp10_81 202000.000000
Rwpos10_82 in10_82 sp10_82 202000.000000
Rwpos10_83 in10_83 sp10_83 202000.000000
Rwpos10_84 in10_84 sp10_84 202000.000000
Rwpos11_1 in11_1 sp11_1 78000.000000
Rwpos11_2 in11_2 sp11_2 78000.000000
Rwpos11_3 in11_3 sp11_3 78000.000000
Rwpos11_4 in11_4 sp11_4 78000.000000
Rwpos11_5 in11_5 sp11_5 78000.000000
Rwpos11_6 in11_6 sp11_6 202000.000000
Rwpos11_7 in11_7 sp11_7 202000.000000
Rwpos11_8 in11_8 sp11_8 78000.000000
Rwpos11_9 in11_9 sp11_9 78000.000000
Rwpos11_10 in11_10 sp11_10 202000.000000
Rwpos11_11 in11_11 sp11_11 202000.000000
Rwpos11_12 in11_12 sp11_12 78000.000000
Rwpos11_13 in11_13 sp11_13 78000.000000
Rwpos11_14 in11_14 sp11_14 202000.000000
Rwpos11_15 in11_15 sp11_15 78000.000000
Rwpos11_16 in11_16 sp11_16 78000.000000
Rwpos11_17 in11_17 sp11_17 202000.000000
Rwpos11_18 in11_18 sp11_18 78000.000000
Rwpos11_19 in11_19 sp11_19 78000.000000
Rwpos11_20 in11_20 sp11_20 78000.000000
Rwpos11_21 in11_21 sp11_21 78000.000000
Rwpos11_22 in11_22 sp11_22 78000.000000
Rwpos11_23 in11_23 sp11_23 78000.000000
Rwpos11_24 in11_24 sp11_24 202000.000000
Rwpos11_25 in11_25 sp11_25 202000.000000
Rwpos11_26 in11_26 sp11_26 78000.000000
Rwpos11_27 in11_27 sp11_27 78000.000000
Rwpos11_28 in11_28 sp11_28 78000.000000
Rwpos11_29 in11_29 sp11_29 202000.000000
Rwpos11_30 in11_30 sp11_30 78000.000000
Rwpos11_31 in11_31 sp11_31 202000.000000
Rwpos11_32 in11_32 sp11_32 78000.000000
Rwpos11_33 in11_33 sp11_33 78000.000000
Rwpos11_34 in11_34 sp11_34 202000.000000
Rwpos11_35 in11_35 sp11_35 78000.000000
Rwpos11_36 in11_36 sp11_36 202000.000000
Rwpos11_37 in11_37 sp11_37 202000.000000
Rwpos11_38 in11_38 sp11_38 78000.000000
Rwpos11_39 in11_39 sp11_39 78000.000000
Rwpos11_40 in11_40 sp11_40 78000.000000
Rwpos11_41 in11_41 sp11_41 78000.000000
Rwpos11_42 in11_42 sp11_42 78000.000000
Rwpos11_43 in11_43 sp11_43 78000.000000
Rwpos11_44 in11_44 sp11_44 202000.000000
Rwpos11_45 in11_45 sp11_45 78000.000000
Rwpos11_46 in11_46 sp11_46 202000.000000
Rwpos11_47 in11_47 sp11_47 78000.000000
Rwpos11_48 in11_48 sp11_48 202000.000000
Rwpos11_49 in11_49 sp11_49 202000.000000
Rwpos11_50 in11_50 sp11_50 202000.000000
Rwpos11_51 in11_51 sp11_51 202000.000000
Rwpos11_52 in11_52 sp11_52 78000.000000
Rwpos11_53 in11_53 sp11_53 202000.000000
Rwpos11_54 in11_54 sp11_54 78000.000000
Rwpos11_55 in11_55 sp11_55 78000.000000
Rwpos11_56 in11_56 sp11_56 202000.000000
Rwpos11_57 in11_57 sp11_57 202000.000000
Rwpos11_58 in11_58 sp11_58 78000.000000
Rwpos11_59 in11_59 sp11_59 202000.000000
Rwpos11_60 in11_60 sp11_60 202000.000000
Rwpos11_61 in11_61 sp11_61 78000.000000
Rwpos11_62 in11_62 sp11_62 202000.000000
Rwpos11_63 in11_63 sp11_63 78000.000000
Rwpos11_64 in11_64 sp11_64 202000.000000
Rwpos11_65 in11_65 sp11_65 202000.000000
Rwpos11_66 in11_66 sp11_66 202000.000000
Rwpos11_67 in11_67 sp11_67 78000.000000
Rwpos11_68 in11_68 sp11_68 78000.000000
Rwpos11_69 in11_69 sp11_69 202000.000000
Rwpos11_70 in11_70 sp11_70 202000.000000
Rwpos11_71 in11_71 sp11_71 202000.000000
Rwpos11_72 in11_72 sp11_72 78000.000000
Rwpos11_73 in11_73 sp11_73 202000.000000
Rwpos11_74 in11_74 sp11_74 78000.000000
Rwpos11_75 in11_75 sp11_75 202000.000000
Rwpos11_76 in11_76 sp11_76 78000.000000
Rwpos11_77 in11_77 sp11_77 78000.000000
Rwpos11_78 in11_78 sp11_78 78000.000000
Rwpos11_79 in11_79 sp11_79 202000.000000
Rwpos11_80 in11_80 sp11_80 78000.000000
Rwpos11_81 in11_81 sp11_81 202000.000000
Rwpos11_82 in11_82 sp11_82 78000.000000
Rwpos11_83 in11_83 sp11_83 78000.000000
Rwpos11_84 in11_84 sp11_84 78000.000000
Rwpos12_1 in12_1 sp12_1 202000.000000
Rwpos12_2 in12_2 sp12_2 202000.000000
Rwpos12_3 in12_3 sp12_3 202000.000000
Rwpos12_4 in12_4 sp12_4 78000.000000
Rwpos12_5 in12_5 sp12_5 202000.000000
Rwpos12_6 in12_6 sp12_6 78000.000000
Rwpos12_7 in12_7 sp12_7 202000.000000
Rwpos12_8 in12_8 sp12_8 78000.000000
Rwpos12_9 in12_9 sp12_9 78000.000000
Rwpos12_10 in12_10 sp12_10 78000.000000
Rwpos12_11 in12_11 sp12_11 78000.000000
Rwpos12_12 in12_12 sp12_12 78000.000000
Rwpos12_13 in12_13 sp12_13 78000.000000
Rwpos12_14 in12_14 sp12_14 202000.000000
Rwpos12_15 in12_15 sp12_15 78000.000000
Rwpos12_16 in12_16 sp12_16 78000.000000
Rwpos12_17 in12_17 sp12_17 202000.000000
Rwpos12_18 in12_18 sp12_18 78000.000000
Rwpos12_19 in12_19 sp12_19 78000.000000
Rwpos12_20 in12_20 sp12_20 78000.000000
Rwpos12_21 in12_21 sp12_21 78000.000000
Rwpos12_22 in12_22 sp12_22 78000.000000
Rwpos12_23 in12_23 sp12_23 78000.000000
Rwpos12_24 in12_24 sp12_24 202000.000000
Rwpos12_25 in12_25 sp12_25 202000.000000
Rwpos12_26 in12_26 sp12_26 202000.000000
Rwpos12_27 in12_27 sp12_27 202000.000000
Rwpos12_28 in12_28 sp12_28 202000.000000
Rwpos12_29 in12_29 sp12_29 78000.000000
Rwpos12_30 in12_30 sp12_30 78000.000000
Rwpos12_31 in12_31 sp12_31 202000.000000
Rwpos12_32 in12_32 sp12_32 202000.000000
Rwpos12_33 in12_33 sp12_33 78000.000000
Rwpos12_34 in12_34 sp12_34 78000.000000
Rwpos12_35 in12_35 sp12_35 202000.000000
Rwpos12_36 in12_36 sp12_36 202000.000000
Rwpos12_37 in12_37 sp12_37 78000.000000
Rwpos12_38 in12_38 sp12_38 78000.000000
Rwpos12_39 in12_39 sp12_39 202000.000000
Rwpos12_40 in12_40 sp12_40 78000.000000
Rwpos12_41 in12_41 sp12_41 202000.000000
Rwpos12_42 in12_42 sp12_42 202000.000000
Rwpos12_43 in12_43 sp12_43 78000.000000
Rwpos12_44 in12_44 sp12_44 202000.000000
Rwpos12_45 in12_45 sp12_45 78000.000000
Rwpos12_46 in12_46 sp12_46 202000.000000
Rwpos12_47 in12_47 sp12_47 202000.000000
Rwpos12_48 in12_48 sp12_48 202000.000000
Rwpos12_49 in12_49 sp12_49 78000.000000
Rwpos12_50 in12_50 sp12_50 202000.000000
Rwpos12_51 in12_51 sp12_51 78000.000000
Rwpos12_52 in12_52 sp12_52 78000.000000
Rwpos12_53 in12_53 sp12_53 202000.000000
Rwpos12_54 in12_54 sp12_54 202000.000000
Rwpos12_55 in12_55 sp12_55 202000.000000
Rwpos12_56 in12_56 sp12_56 78000.000000
Rwpos12_57 in12_57 sp12_57 78000.000000
Rwpos12_58 in12_58 sp12_58 78000.000000
Rwpos12_59 in12_59 sp12_59 78000.000000
Rwpos12_60 in12_60 sp12_60 202000.000000
Rwpos12_61 in12_61 sp12_61 78000.000000
Rwpos12_62 in12_62 sp12_62 202000.000000
Rwpos12_63 in12_63 sp12_63 78000.000000
Rwpos12_64 in12_64 sp12_64 78000.000000
Rwpos12_65 in12_65 sp12_65 202000.000000
Rwpos12_66 in12_66 sp12_66 78000.000000
Rwpos12_67 in12_67 sp12_67 202000.000000
Rwpos12_68 in12_68 sp12_68 78000.000000
Rwpos12_69 in12_69 sp12_69 78000.000000
Rwpos12_70 in12_70 sp12_70 78000.000000
Rwpos12_71 in12_71 sp12_71 78000.000000
Rwpos12_72 in12_72 sp12_72 202000.000000
Rwpos12_73 in12_73 sp12_73 78000.000000
Rwpos12_74 in12_74 sp12_74 202000.000000
Rwpos12_75 in12_75 sp12_75 202000.000000
Rwpos12_76 in12_76 sp12_76 202000.000000
Rwpos12_77 in12_77 sp12_77 78000.000000
Rwpos12_78 in12_78 sp12_78 78000.000000
Rwpos12_79 in12_79 sp12_79 78000.000000
Rwpos12_80 in12_80 sp12_80 78000.000000
Rwpos12_81 in12_81 sp12_81 202000.000000
Rwpos12_82 in12_82 sp12_82 78000.000000
Rwpos12_83 in12_83 sp12_83 78000.000000
Rwpos12_84 in12_84 sp12_84 78000.000000
Rwpos13_1 in13_1 sp13_1 78000.000000
Rwpos13_2 in13_2 sp13_2 78000.000000
Rwpos13_3 in13_3 sp13_3 202000.000000
Rwpos13_4 in13_4 sp13_4 78000.000000
Rwpos13_5 in13_5 sp13_5 78000.000000
Rwpos13_6 in13_6 sp13_6 202000.000000
Rwpos13_7 in13_7 sp13_7 78000.000000
Rwpos13_8 in13_8 sp13_8 78000.000000
Rwpos13_9 in13_9 sp13_9 78000.000000
Rwpos13_10 in13_10 sp13_10 202000.000000
Rwpos13_11 in13_11 sp13_11 202000.000000
Rwpos13_12 in13_12 sp13_12 78000.000000
Rwpos13_13 in13_13 sp13_13 202000.000000
Rwpos13_14 in13_14 sp13_14 202000.000000
Rwpos13_15 in13_15 sp13_15 202000.000000
Rwpos13_16 in13_16 sp13_16 78000.000000
Rwpos13_17 in13_17 sp13_17 202000.000000
Rwpos13_18 in13_18 sp13_18 78000.000000
Rwpos13_19 in13_19 sp13_19 202000.000000
Rwpos13_20 in13_20 sp13_20 202000.000000
Rwpos13_21 in13_21 sp13_21 78000.000000
Rwpos13_22 in13_22 sp13_22 78000.000000
Rwpos13_23 in13_23 sp13_23 202000.000000
Rwpos13_24 in13_24 sp13_24 202000.000000
Rwpos13_25 in13_25 sp13_25 78000.000000
Rwpos13_26 in13_26 sp13_26 202000.000000
Rwpos13_27 in13_27 sp13_27 78000.000000
Rwpos13_28 in13_28 sp13_28 202000.000000
Rwpos13_29 in13_29 sp13_29 78000.000000
Rwpos13_30 in13_30 sp13_30 78000.000000
Rwpos13_31 in13_31 sp13_31 78000.000000
Rwpos13_32 in13_32 sp13_32 202000.000000
Rwpos13_33 in13_33 sp13_33 202000.000000
Rwpos13_34 in13_34 sp13_34 202000.000000
Rwpos13_35 in13_35 sp13_35 78000.000000
Rwpos13_36 in13_36 sp13_36 78000.000000
Rwpos13_37 in13_37 sp13_37 78000.000000
Rwpos13_38 in13_38 sp13_38 202000.000000
Rwpos13_39 in13_39 sp13_39 202000.000000
Rwpos13_40 in13_40 sp13_40 202000.000000
Rwpos13_41 in13_41 sp13_41 78000.000000
Rwpos13_42 in13_42 sp13_42 78000.000000
Rwpos13_43 in13_43 sp13_43 78000.000000
Rwpos13_44 in13_44 sp13_44 78000.000000
Rwpos13_45 in13_45 sp13_45 202000.000000
Rwpos13_46 in13_46 sp13_46 202000.000000
Rwpos13_47 in13_47 sp13_47 202000.000000
Rwpos13_48 in13_48 sp13_48 202000.000000
Rwpos13_49 in13_49 sp13_49 78000.000000
Rwpos13_50 in13_50 sp13_50 202000.000000
Rwpos13_51 in13_51 sp13_51 78000.000000
Rwpos13_52 in13_52 sp13_52 78000.000000
Rwpos13_53 in13_53 sp13_53 78000.000000
Rwpos13_54 in13_54 sp13_54 78000.000000
Rwpos13_55 in13_55 sp13_55 202000.000000
Rwpos13_56 in13_56 sp13_56 78000.000000
Rwpos13_57 in13_57 sp13_57 78000.000000
Rwpos13_58 in13_58 sp13_58 202000.000000
Rwpos13_59 in13_59 sp13_59 78000.000000
Rwpos13_60 in13_60 sp13_60 78000.000000
Rwpos13_61 in13_61 sp13_61 78000.000000
Rwpos13_62 in13_62 sp13_62 78000.000000
Rwpos13_63 in13_63 sp13_63 78000.000000
Rwpos13_64 in13_64 sp13_64 78000.000000
Rwpos13_65 in13_65 sp13_65 78000.000000
Rwpos13_66 in13_66 sp13_66 78000.000000
Rwpos13_67 in13_67 sp13_67 202000.000000
Rwpos13_68 in13_68 sp13_68 78000.000000
Rwpos13_69 in13_69 sp13_69 78000.000000
Rwpos13_70 in13_70 sp13_70 78000.000000
Rwpos13_71 in13_71 sp13_71 78000.000000
Rwpos13_72 in13_72 sp13_72 78000.000000
Rwpos13_73 in13_73 sp13_73 78000.000000
Rwpos13_74 in13_74 sp13_74 202000.000000
Rwpos13_75 in13_75 sp13_75 202000.000000
Rwpos13_76 in13_76 sp13_76 78000.000000
Rwpos13_77 in13_77 sp13_77 202000.000000
Rwpos13_78 in13_78 sp13_78 78000.000000
Rwpos13_79 in13_79 sp13_79 78000.000000
Rwpos13_80 in13_80 sp13_80 78000.000000
Rwpos13_81 in13_81 sp13_81 202000.000000
Rwpos13_82 in13_82 sp13_82 78000.000000
Rwpos13_83 in13_83 sp13_83 202000.000000
Rwpos13_84 in13_84 sp13_84 78000.000000
Rwpos14_1 in14_1 sp14_1 78000.000000
Rwpos14_2 in14_2 sp14_2 78000.000000
Rwpos14_3 in14_3 sp14_3 78000.000000
Rwpos14_4 in14_4 sp14_4 202000.000000
Rwpos14_5 in14_5 sp14_5 202000.000000
Rwpos14_6 in14_6 sp14_6 78000.000000
Rwpos14_7 in14_7 sp14_7 78000.000000
Rwpos14_8 in14_8 sp14_8 202000.000000
Rwpos14_9 in14_9 sp14_9 202000.000000
Rwpos14_10 in14_10 sp14_10 202000.000000
Rwpos14_11 in14_11 sp14_11 78000.000000
Rwpos14_12 in14_12 sp14_12 202000.000000
Rwpos14_13 in14_13 sp14_13 202000.000000
Rwpos14_14 in14_14 sp14_14 78000.000000
Rwpos14_15 in14_15 sp14_15 202000.000000
Rwpos14_16 in14_16 sp14_16 78000.000000
Rwpos14_17 in14_17 sp14_17 78000.000000
Rwpos14_18 in14_18 sp14_18 202000.000000
Rwpos14_19 in14_19 sp14_19 78000.000000
Rwpos14_20 in14_20 sp14_20 202000.000000
Rwpos14_21 in14_21 sp14_21 78000.000000
Rwpos14_22 in14_22 sp14_22 78000.000000
Rwpos14_23 in14_23 sp14_23 78000.000000
Rwpos14_24 in14_24 sp14_24 202000.000000
Rwpos14_25 in14_25 sp14_25 78000.000000
Rwpos14_26 in14_26 sp14_26 78000.000000
Rwpos14_27 in14_27 sp14_27 202000.000000
Rwpos14_28 in14_28 sp14_28 202000.000000
Rwpos14_29 in14_29 sp14_29 78000.000000
Rwpos14_30 in14_30 sp14_30 78000.000000
Rwpos14_31 in14_31 sp14_31 78000.000000
Rwpos14_32 in14_32 sp14_32 202000.000000
Rwpos14_33 in14_33 sp14_33 78000.000000
Rwpos14_34 in14_34 sp14_34 78000.000000
Rwpos14_35 in14_35 sp14_35 202000.000000
Rwpos14_36 in14_36 sp14_36 202000.000000
Rwpos14_37 in14_37 sp14_37 78000.000000
Rwpos14_38 in14_38 sp14_38 78000.000000
Rwpos14_39 in14_39 sp14_39 202000.000000
Rwpos14_40 in14_40 sp14_40 78000.000000
Rwpos14_41 in14_41 sp14_41 202000.000000
Rwpos14_42 in14_42 sp14_42 78000.000000
Rwpos14_43 in14_43 sp14_43 78000.000000
Rwpos14_44 in14_44 sp14_44 78000.000000
Rwpos14_45 in14_45 sp14_45 202000.000000
Rwpos14_46 in14_46 sp14_46 78000.000000
Rwpos14_47 in14_47 sp14_47 78000.000000
Rwpos14_48 in14_48 sp14_48 202000.000000
Rwpos14_49 in14_49 sp14_49 78000.000000
Rwpos14_50 in14_50 sp14_50 78000.000000
Rwpos14_51 in14_51 sp14_51 78000.000000
Rwpos14_52 in14_52 sp14_52 78000.000000
Rwpos14_53 in14_53 sp14_53 78000.000000
Rwpos14_54 in14_54 sp14_54 202000.000000
Rwpos14_55 in14_55 sp14_55 78000.000000
Rwpos14_56 in14_56 sp14_56 202000.000000
Rwpos14_57 in14_57 sp14_57 78000.000000
Rwpos14_58 in14_58 sp14_58 78000.000000
Rwpos14_59 in14_59 sp14_59 78000.000000
Rwpos14_60 in14_60 sp14_60 202000.000000
Rwpos14_61 in14_61 sp14_61 78000.000000
Rwpos14_62 in14_62 sp14_62 78000.000000
Rwpos14_63 in14_63 sp14_63 202000.000000
Rwpos14_64 in14_64 sp14_64 78000.000000
Rwpos14_65 in14_65 sp14_65 202000.000000
Rwpos14_66 in14_66 sp14_66 78000.000000
Rwpos14_67 in14_67 sp14_67 202000.000000
Rwpos14_68 in14_68 sp14_68 202000.000000
Rwpos14_69 in14_69 sp14_69 202000.000000
Rwpos14_70 in14_70 sp14_70 202000.000000
Rwpos14_71 in14_71 sp14_71 202000.000000
Rwpos14_72 in14_72 sp14_72 78000.000000
Rwpos14_73 in14_73 sp14_73 78000.000000
Rwpos14_74 in14_74 sp14_74 78000.000000
Rwpos14_75 in14_75 sp14_75 202000.000000
Rwpos14_76 in14_76 sp14_76 78000.000000
Rwpos14_77 in14_77 sp14_77 78000.000000
Rwpos14_78 in14_78 sp14_78 78000.000000
Rwpos14_79 in14_79 sp14_79 202000.000000
Rwpos14_80 in14_80 sp14_80 202000.000000
Rwpos14_81 in14_81 sp14_81 202000.000000
Rwpos14_82 in14_82 sp14_82 202000.000000
Rwpos14_83 in14_83 sp14_83 78000.000000
Rwpos14_84 in14_84 sp14_84 202000.000000
Rwpos15_1 in15_1 sp15_1 78000.000000
Rwpos15_2 in15_2 sp15_2 78000.000000
Rwpos15_3 in15_3 sp15_3 78000.000000
Rwpos15_4 in15_4 sp15_4 202000.000000
Rwpos15_5 in15_5 sp15_5 202000.000000
Rwpos15_6 in15_6 sp15_6 78000.000000
Rwpos15_7 in15_7 sp15_7 78000.000000
Rwpos15_8 in15_8 sp15_8 202000.000000
Rwpos15_9 in15_9 sp15_9 202000.000000
Rwpos15_10 in15_10 sp15_10 202000.000000
Rwpos15_11 in15_11 sp15_11 78000.000000
Rwpos15_12 in15_12 sp15_12 78000.000000
Rwpos15_13 in15_13 sp15_13 202000.000000
Rwpos15_14 in15_14 sp15_14 202000.000000
Rwpos15_15 in15_15 sp15_15 78000.000000
Rwpos15_16 in15_16 sp15_16 78000.000000
Rwpos15_17 in15_17 sp15_17 78000.000000
Rwpos15_18 in15_18 sp15_18 202000.000000
Rwpos15_19 in15_19 sp15_19 78000.000000
Rwpos15_20 in15_20 sp15_20 202000.000000
Rwpos15_21 in15_21 sp15_21 78000.000000
Rwpos15_22 in15_22 sp15_22 78000.000000
Rwpos15_23 in15_23 sp15_23 202000.000000
Rwpos15_24 in15_24 sp15_24 78000.000000
Rwpos15_25 in15_25 sp15_25 78000.000000
Rwpos15_26 in15_26 sp15_26 202000.000000
Rwpos15_27 in15_27 sp15_27 202000.000000
Rwpos15_28 in15_28 sp15_28 78000.000000
Rwpos15_29 in15_29 sp15_29 78000.000000
Rwpos15_30 in15_30 sp15_30 202000.000000
Rwpos15_31 in15_31 sp15_31 202000.000000
Rwpos15_32 in15_32 sp15_32 202000.000000
Rwpos15_33 in15_33 sp15_33 78000.000000
Rwpos15_34 in15_34 sp15_34 78000.000000
Rwpos15_35 in15_35 sp15_35 78000.000000
Rwpos15_36 in15_36 sp15_36 78000.000000
Rwpos15_37 in15_37 sp15_37 78000.000000
Rwpos15_38 in15_38 sp15_38 202000.000000
Rwpos15_39 in15_39 sp15_39 202000.000000
Rwpos15_40 in15_40 sp15_40 78000.000000
Rwpos15_41 in15_41 sp15_41 202000.000000
Rwpos15_42 in15_42 sp15_42 78000.000000
Rwpos15_43 in15_43 sp15_43 78000.000000
Rwpos15_44 in15_44 sp15_44 78000.000000
Rwpos15_45 in15_45 sp15_45 78000.000000
Rwpos15_46 in15_46 sp15_46 202000.000000
Rwpos15_47 in15_47 sp15_47 78000.000000
Rwpos15_48 in15_48 sp15_48 202000.000000
Rwpos15_49 in15_49 sp15_49 78000.000000
Rwpos15_50 in15_50 sp15_50 202000.000000
Rwpos15_51 in15_51 sp15_51 78000.000000
Rwpos15_52 in15_52 sp15_52 78000.000000
Rwpos15_53 in15_53 sp15_53 202000.000000
Rwpos15_54 in15_54 sp15_54 202000.000000
Rwpos15_55 in15_55 sp15_55 202000.000000
Rwpos15_56 in15_56 sp15_56 78000.000000
Rwpos15_57 in15_57 sp15_57 78000.000000
Rwpos15_58 in15_58 sp15_58 78000.000000
Rwpos15_59 in15_59 sp15_59 202000.000000
Rwpos15_60 in15_60 sp15_60 78000.000000
Rwpos15_61 in15_61 sp15_61 78000.000000
Rwpos15_62 in15_62 sp15_62 202000.000000
Rwpos15_63 in15_63 sp15_63 78000.000000
Rwpos15_64 in15_64 sp15_64 202000.000000
Rwpos15_65 in15_65 sp15_65 202000.000000
Rwpos15_66 in15_66 sp15_66 78000.000000
Rwpos15_67 in15_67 sp15_67 78000.000000
Rwpos15_68 in15_68 sp15_68 78000.000000
Rwpos15_69 in15_69 sp15_69 78000.000000
Rwpos15_70 in15_70 sp15_70 78000.000000
Rwpos15_71 in15_71 sp15_71 78000.000000
Rwpos15_72 in15_72 sp15_72 78000.000000
Rwpos15_73 in15_73 sp15_73 78000.000000
Rwpos15_74 in15_74 sp15_74 78000.000000
Rwpos15_75 in15_75 sp15_75 78000.000000
Rwpos15_76 in15_76 sp15_76 78000.000000
Rwpos15_77 in15_77 sp15_77 202000.000000
Rwpos15_78 in15_78 sp15_78 78000.000000
Rwpos15_79 in15_79 sp15_79 78000.000000
Rwpos15_80 in15_80 sp15_80 202000.000000
Rwpos15_81 in15_81 sp15_81 78000.000000
Rwpos15_82 in15_82 sp15_82 202000.000000
Rwpos15_83 in15_83 sp15_83 78000.000000
Rwpos15_84 in15_84 sp15_84 202000.000000
Rwpos16_1 in16_1 sp16_1 202000.000000
Rwpos16_2 in16_2 sp16_2 202000.000000
Rwpos16_3 in16_3 sp16_3 202000.000000
Rwpos16_4 in16_4 sp16_4 78000.000000
Rwpos16_5 in16_5 sp16_5 78000.000000
Rwpos16_6 in16_6 sp16_6 78000.000000
Rwpos16_7 in16_7 sp16_7 78000.000000
Rwpos16_8 in16_8 sp16_8 202000.000000
Rwpos16_9 in16_9 sp16_9 202000.000000
Rwpos16_10 in16_10 sp16_10 78000.000000
Rwpos16_11 in16_11 sp16_11 78000.000000
Rwpos16_12 in16_12 sp16_12 78000.000000
Rwpos16_13 in16_13 sp16_13 202000.000000
Rwpos16_14 in16_14 sp16_14 78000.000000
Rwpos16_15 in16_15 sp16_15 78000.000000
Rwpos16_16 in16_16 sp16_16 78000.000000
Rwpos16_17 in16_17 sp16_17 78000.000000
Rwpos16_18 in16_18 sp16_18 202000.000000
Rwpos16_19 in16_19 sp16_19 78000.000000
Rwpos16_20 in16_20 sp16_20 78000.000000
Rwpos16_21 in16_21 sp16_21 78000.000000
Rwpos16_22 in16_22 sp16_22 78000.000000
Rwpos16_23 in16_23 sp16_23 78000.000000
Rwpos16_24 in16_24 sp16_24 202000.000000
Rwpos16_25 in16_25 sp16_25 78000.000000
Rwpos16_26 in16_26 sp16_26 202000.000000
Rwpos16_27 in16_27 sp16_27 78000.000000
Rwpos16_28 in16_28 sp16_28 78000.000000
Rwpos16_29 in16_29 sp16_29 202000.000000
Rwpos16_30 in16_30 sp16_30 78000.000000
Rwpos16_31 in16_31 sp16_31 78000.000000
Rwpos16_32 in16_32 sp16_32 78000.000000
Rwpos16_33 in16_33 sp16_33 202000.000000
Rwpos16_34 in16_34 sp16_34 78000.000000
Rwpos16_35 in16_35 sp16_35 202000.000000
Rwpos16_36 in16_36 sp16_36 202000.000000
Rwpos16_37 in16_37 sp16_37 78000.000000
Rwpos16_38 in16_38 sp16_38 78000.000000
Rwpos16_39 in16_39 sp16_39 202000.000000
Rwpos16_40 in16_40 sp16_40 78000.000000
Rwpos16_41 in16_41 sp16_41 78000.000000
Rwpos16_42 in16_42 sp16_42 202000.000000
Rwpos16_43 in16_43 sp16_43 78000.000000
Rwpos16_44 in16_44 sp16_44 78000.000000
Rwpos16_45 in16_45 sp16_45 78000.000000
Rwpos16_46 in16_46 sp16_46 78000.000000
Rwpos16_47 in16_47 sp16_47 202000.000000
Rwpos16_48 in16_48 sp16_48 78000.000000
Rwpos16_49 in16_49 sp16_49 202000.000000
Rwpos16_50 in16_50 sp16_50 78000.000000
Rwpos16_51 in16_51 sp16_51 78000.000000
Rwpos16_52 in16_52 sp16_52 202000.000000
Rwpos16_53 in16_53 sp16_53 202000.000000
Rwpos16_54 in16_54 sp16_54 78000.000000
Rwpos16_55 in16_55 sp16_55 202000.000000
Rwpos16_56 in16_56 sp16_56 78000.000000
Rwpos16_57 in16_57 sp16_57 78000.000000
Rwpos16_58 in16_58 sp16_58 78000.000000
Rwpos16_59 in16_59 sp16_59 78000.000000
Rwpos16_60 in16_60 sp16_60 202000.000000
Rwpos16_61 in16_61 sp16_61 202000.000000
Rwpos16_62 in16_62 sp16_62 78000.000000
Rwpos16_63 in16_63 sp16_63 202000.000000
Rwpos16_64 in16_64 sp16_64 202000.000000
Rwpos16_65 in16_65 sp16_65 78000.000000
Rwpos16_66 in16_66 sp16_66 202000.000000
Rwpos16_67 in16_67 sp16_67 202000.000000
Rwpos16_68 in16_68 sp16_68 78000.000000
Rwpos16_69 in16_69 sp16_69 78000.000000
Rwpos16_70 in16_70 sp16_70 78000.000000
Rwpos16_71 in16_71 sp16_71 78000.000000
Rwpos16_72 in16_72 sp16_72 78000.000000
Rwpos16_73 in16_73 sp16_73 78000.000000
Rwpos16_74 in16_74 sp16_74 202000.000000
Rwpos16_75 in16_75 sp16_75 78000.000000
Rwpos16_76 in16_76 sp16_76 202000.000000
Rwpos16_77 in16_77 sp16_77 78000.000000
Rwpos16_78 in16_78 sp16_78 78000.000000
Rwpos16_79 in16_79 sp16_79 78000.000000
Rwpos16_80 in16_80 sp16_80 202000.000000
Rwpos16_81 in16_81 sp16_81 78000.000000
Rwpos16_82 in16_82 sp16_82 202000.000000
Rwpos16_83 in16_83 sp16_83 202000.000000
Rwpos16_84 in16_84 sp16_84 78000.000000
Rwpos17_1 in17_1 sp17_1 78000.000000
Rwpos17_2 in17_2 sp17_2 78000.000000
Rwpos17_3 in17_3 sp17_3 202000.000000
Rwpos17_4 in17_4 sp17_4 78000.000000
Rwpos17_5 in17_5 sp17_5 78000.000000
Rwpos17_6 in17_6 sp17_6 78000.000000
Rwpos17_7 in17_7 sp17_7 202000.000000
Rwpos17_8 in17_8 sp17_8 78000.000000
Rwpos17_9 in17_9 sp17_9 78000.000000
Rwpos17_10 in17_10 sp17_10 78000.000000
Rwpos17_11 in17_11 sp17_11 202000.000000
Rwpos17_12 in17_12 sp17_12 78000.000000
Rwpos17_13 in17_13 sp17_13 78000.000000
Rwpos17_14 in17_14 sp17_14 202000.000000
Rwpos17_15 in17_15 sp17_15 202000.000000
Rwpos17_16 in17_16 sp17_16 78000.000000
Rwpos17_17 in17_17 sp17_17 202000.000000
Rwpos17_18 in17_18 sp17_18 78000.000000
Rwpos17_19 in17_19 sp17_19 78000.000000
Rwpos17_20 in17_20 sp17_20 78000.000000
Rwpos17_21 in17_21 sp17_21 78000.000000
Rwpos17_22 in17_22 sp17_22 78000.000000
Rwpos17_23 in17_23 sp17_23 78000.000000
Rwpos17_24 in17_24 sp17_24 202000.000000
Rwpos17_25 in17_25 sp17_25 202000.000000
Rwpos17_26 in17_26 sp17_26 78000.000000
Rwpos17_27 in17_27 sp17_27 78000.000000
Rwpos17_28 in17_28 sp17_28 78000.000000
Rwpos17_29 in17_29 sp17_29 78000.000000
Rwpos17_30 in17_30 sp17_30 202000.000000
Rwpos17_31 in17_31 sp17_31 202000.000000
Rwpos17_32 in17_32 sp17_32 78000.000000
Rwpos17_33 in17_33 sp17_33 202000.000000
Rwpos17_34 in17_34 sp17_34 78000.000000
Rwpos17_35 in17_35 sp17_35 202000.000000
Rwpos17_36 in17_36 sp17_36 78000.000000
Rwpos17_37 in17_37 sp17_37 78000.000000
Rwpos17_38 in17_38 sp17_38 78000.000000
Rwpos17_39 in17_39 sp17_39 78000.000000
Rwpos17_40 in17_40 sp17_40 78000.000000
Rwpos17_41 in17_41 sp17_41 78000.000000
Rwpos17_42 in17_42 sp17_42 78000.000000
Rwpos17_43 in17_43 sp17_43 202000.000000
Rwpos17_44 in17_44 sp17_44 78000.000000
Rwpos17_45 in17_45 sp17_45 78000.000000
Rwpos17_46 in17_46 sp17_46 202000.000000
Rwpos17_47 in17_47 sp17_47 202000.000000
Rwpos17_48 in17_48 sp17_48 78000.000000
Rwpos17_49 in17_49 sp17_49 202000.000000
Rwpos17_50 in17_50 sp17_50 202000.000000
Rwpos17_51 in17_51 sp17_51 202000.000000
Rwpos17_52 in17_52 sp17_52 202000.000000
Rwpos17_53 in17_53 sp17_53 202000.000000
Rwpos17_54 in17_54 sp17_54 202000.000000
Rwpos17_55 in17_55 sp17_55 78000.000000
Rwpos17_56 in17_56 sp17_56 78000.000000
Rwpos17_57 in17_57 sp17_57 202000.000000
Rwpos17_58 in17_58 sp17_58 78000.000000
Rwpos17_59 in17_59 sp17_59 202000.000000
Rwpos17_60 in17_60 sp17_60 78000.000000
Rwpos17_61 in17_61 sp17_61 78000.000000
Rwpos17_62 in17_62 sp17_62 202000.000000
Rwpos17_63 in17_63 sp17_63 78000.000000
Rwpos17_64 in17_64 sp17_64 78000.000000
Rwpos17_65 in17_65 sp17_65 78000.000000
Rwpos17_66 in17_66 sp17_66 78000.000000
Rwpos17_67 in17_67 sp17_67 202000.000000
Rwpos17_68 in17_68 sp17_68 78000.000000
Rwpos17_69 in17_69 sp17_69 202000.000000
Rwpos17_70 in17_70 sp17_70 78000.000000
Rwpos17_71 in17_71 sp17_71 78000.000000
Rwpos17_72 in17_72 sp17_72 202000.000000
Rwpos17_73 in17_73 sp17_73 78000.000000
Rwpos17_74 in17_74 sp17_74 202000.000000
Rwpos17_75 in17_75 sp17_75 202000.000000
Rwpos17_76 in17_76 sp17_76 202000.000000
Rwpos17_77 in17_77 sp17_77 78000.000000
Rwpos17_78 in17_78 sp17_78 78000.000000
Rwpos17_79 in17_79 sp17_79 78000.000000
Rwpos17_80 in17_80 sp17_80 78000.000000
Rwpos17_81 in17_81 sp17_81 202000.000000
Rwpos17_82 in17_82 sp17_82 78000.000000
Rwpos17_83 in17_83 sp17_83 78000.000000
Rwpos17_84 in17_84 sp17_84 78000.000000
Rwpos18_1 in18_1 sp18_1 202000.000000
Rwpos18_2 in18_2 sp18_2 78000.000000
Rwpos18_3 in18_3 sp18_3 78000.000000
Rwpos18_4 in18_4 sp18_4 202000.000000
Rwpos18_5 in18_5 sp18_5 202000.000000
Rwpos18_6 in18_6 sp18_6 202000.000000
Rwpos18_7 in18_7 sp18_7 78000.000000
Rwpos18_8 in18_8 sp18_8 78000.000000
Rwpos18_9 in18_9 sp18_9 202000.000000
Rwpos18_10 in18_10 sp18_10 78000.000000
Rwpos18_11 in18_11 sp18_11 78000.000000
Rwpos18_12 in18_12 sp18_12 202000.000000
Rwpos18_13 in18_13 sp18_13 202000.000000
Rwpos18_14 in18_14 sp18_14 202000.000000
Rwpos18_15 in18_15 sp18_15 202000.000000
Rwpos18_16 in18_16 sp18_16 202000.000000
Rwpos18_17 in18_17 sp18_17 202000.000000
Rwpos18_18 in18_18 sp18_18 202000.000000
Rwpos18_19 in18_19 sp18_19 202000.000000
Rwpos18_20 in18_20 sp18_20 202000.000000
Rwpos18_21 in18_21 sp18_21 78000.000000
Rwpos18_22 in18_22 sp18_22 202000.000000
Rwpos18_23 in18_23 sp18_23 78000.000000
Rwpos18_24 in18_24 sp18_24 202000.000000
Rwpos18_25 in18_25 sp18_25 78000.000000
Rwpos18_26 in18_26 sp18_26 202000.000000
Rwpos18_27 in18_27 sp18_27 202000.000000
Rwpos18_28 in18_28 sp18_28 202000.000000
Rwpos18_29 in18_29 sp18_29 202000.000000
Rwpos18_30 in18_30 sp18_30 202000.000000
Rwpos18_31 in18_31 sp18_31 202000.000000
Rwpos18_32 in18_32 sp18_32 202000.000000
Rwpos18_33 in18_33 sp18_33 78000.000000
Rwpos18_34 in18_34 sp18_34 202000.000000
Rwpos18_35 in18_35 sp18_35 202000.000000
Rwpos18_36 in18_36 sp18_36 202000.000000
Rwpos18_37 in18_37 sp18_37 78000.000000
Rwpos18_38 in18_38 sp18_38 202000.000000
Rwpos18_39 in18_39 sp18_39 202000.000000
Rwpos18_40 in18_40 sp18_40 78000.000000
Rwpos18_41 in18_41 sp18_41 78000.000000
Rwpos18_42 in18_42 sp18_42 78000.000000
Rwpos18_43 in18_43 sp18_43 78000.000000
Rwpos18_44 in18_44 sp18_44 78000.000000
Rwpos18_45 in18_45 sp18_45 202000.000000
Rwpos18_46 in18_46 sp18_46 78000.000000
Rwpos18_47 in18_47 sp18_47 202000.000000
Rwpos18_48 in18_48 sp18_48 202000.000000
Rwpos18_49 in18_49 sp18_49 78000.000000
Rwpos18_50 in18_50 sp18_50 78000.000000
Rwpos18_51 in18_51 sp18_51 78000.000000
Rwpos18_52 in18_52 sp18_52 78000.000000
Rwpos18_53 in18_53 sp18_53 78000.000000
Rwpos18_54 in18_54 sp18_54 202000.000000
Rwpos18_55 in18_55 sp18_55 202000.000000
Rwpos18_56 in18_56 sp18_56 202000.000000
Rwpos18_57 in18_57 sp18_57 202000.000000
Rwpos18_58 in18_58 sp18_58 78000.000000
Rwpos18_59 in18_59 sp18_59 202000.000000
Rwpos18_60 in18_60 sp18_60 78000.000000
Rwpos18_61 in18_61 sp18_61 78000.000000
Rwpos18_62 in18_62 sp18_62 202000.000000
Rwpos18_63 in18_63 sp18_63 78000.000000
Rwpos18_64 in18_64 sp18_64 202000.000000
Rwpos18_65 in18_65 sp18_65 202000.000000
Rwpos18_66 in18_66 sp18_66 78000.000000
Rwpos18_67 in18_67 sp18_67 202000.000000
Rwpos18_68 in18_68 sp18_68 202000.000000
Rwpos18_69 in18_69 sp18_69 202000.000000
Rwpos18_70 in18_70 sp18_70 78000.000000
Rwpos18_71 in18_71 sp18_71 202000.000000
Rwpos18_72 in18_72 sp18_72 202000.000000
Rwpos18_73 in18_73 sp18_73 78000.000000
Rwpos18_74 in18_74 sp18_74 78000.000000
Rwpos18_75 in18_75 sp18_75 202000.000000
Rwpos18_76 in18_76 sp18_76 78000.000000
Rwpos18_77 in18_77 sp18_77 202000.000000
Rwpos18_78 in18_78 sp18_78 78000.000000
Rwpos18_79 in18_79 sp18_79 78000.000000
Rwpos18_80 in18_80 sp18_80 202000.000000
Rwpos18_81 in18_81 sp18_81 78000.000000
Rwpos18_82 in18_82 sp18_82 202000.000000
Rwpos18_83 in18_83 sp18_83 78000.000000
Rwpos18_84 in18_84 sp18_84 78000.000000
Rwpos19_1 in19_1 sp19_1 78000.000000
Rwpos19_2 in19_2 sp19_2 78000.000000
Rwpos19_3 in19_3 sp19_3 78000.000000
Rwpos19_4 in19_4 sp19_4 78000.000000
Rwpos19_5 in19_5 sp19_5 202000.000000
Rwpos19_6 in19_6 sp19_6 202000.000000
Rwpos19_7 in19_7 sp19_7 202000.000000
Rwpos19_8 in19_8 sp19_8 78000.000000
Rwpos19_9 in19_9 sp19_9 78000.000000
Rwpos19_10 in19_10 sp19_10 78000.000000
Rwpos19_11 in19_11 sp19_11 78000.000000
Rwpos19_12 in19_12 sp19_12 202000.000000
Rwpos19_13 in19_13 sp19_13 78000.000000
Rwpos19_14 in19_14 sp19_14 78000.000000
Rwpos19_15 in19_15 sp19_15 78000.000000
Rwpos19_16 in19_16 sp19_16 202000.000000
Rwpos19_17 in19_17 sp19_17 202000.000000
Rwpos19_18 in19_18 sp19_18 78000.000000
Rwpos19_19 in19_19 sp19_19 202000.000000
Rwpos19_20 in19_20 sp19_20 78000.000000
Rwpos19_21 in19_21 sp19_21 202000.000000
Rwpos19_22 in19_22 sp19_22 78000.000000
Rwpos19_23 in19_23 sp19_23 202000.000000
Rwpos19_24 in19_24 sp19_24 202000.000000
Rwpos19_25 in19_25 sp19_25 78000.000000
Rwpos19_26 in19_26 sp19_26 78000.000000
Rwpos19_27 in19_27 sp19_27 78000.000000
Rwpos19_28 in19_28 sp19_28 202000.000000
Rwpos19_29 in19_29 sp19_29 78000.000000
Rwpos19_30 in19_30 sp19_30 202000.000000
Rwpos19_31 in19_31 sp19_31 202000.000000
Rwpos19_32 in19_32 sp19_32 202000.000000
Rwpos19_33 in19_33 sp19_33 78000.000000
Rwpos19_34 in19_34 sp19_34 202000.000000
Rwpos19_35 in19_35 sp19_35 78000.000000
Rwpos19_36 in19_36 sp19_36 78000.000000
Rwpos19_37 in19_37 sp19_37 202000.000000
Rwpos19_38 in19_38 sp19_38 202000.000000
Rwpos19_39 in19_39 sp19_39 78000.000000
Rwpos19_40 in19_40 sp19_40 202000.000000
Rwpos19_41 in19_41 sp19_41 202000.000000
Rwpos19_42 in19_42 sp19_42 78000.000000
Rwpos19_43 in19_43 sp19_43 78000.000000
Rwpos19_44 in19_44 sp19_44 202000.000000
Rwpos19_45 in19_45 sp19_45 78000.000000
Rwpos19_46 in19_46 sp19_46 78000.000000
Rwpos19_47 in19_47 sp19_47 202000.000000
Rwpos19_48 in19_48 sp19_48 202000.000000
Rwpos19_49 in19_49 sp19_49 78000.000000
Rwpos19_50 in19_50 sp19_50 202000.000000
Rwpos19_51 in19_51 sp19_51 202000.000000
Rwpos19_52 in19_52 sp19_52 202000.000000
Rwpos19_53 in19_53 sp19_53 202000.000000
Rwpos19_54 in19_54 sp19_54 202000.000000
Rwpos19_55 in19_55 sp19_55 202000.000000
Rwpos19_56 in19_56 sp19_56 78000.000000
Rwpos19_57 in19_57 sp19_57 78000.000000
Rwpos19_58 in19_58 sp19_58 202000.000000
Rwpos19_59 in19_59 sp19_59 78000.000000
Rwpos19_60 in19_60 sp19_60 78000.000000
Rwpos19_61 in19_61 sp19_61 78000.000000
Rwpos19_62 in19_62 sp19_62 202000.000000
Rwpos19_63 in19_63 sp19_63 78000.000000
Rwpos19_64 in19_64 sp19_64 78000.000000
Rwpos19_65 in19_65 sp19_65 78000.000000
Rwpos19_66 in19_66 sp19_66 78000.000000
Rwpos19_67 in19_67 sp19_67 202000.000000
Rwpos19_68 in19_68 sp19_68 202000.000000
Rwpos19_69 in19_69 sp19_69 78000.000000
Rwpos19_70 in19_70 sp19_70 78000.000000
Rwpos19_71 in19_71 sp19_71 78000.000000
Rwpos19_72 in19_72 sp19_72 202000.000000
Rwpos19_73 in19_73 sp19_73 202000.000000
Rwpos19_74 in19_74 sp19_74 78000.000000
Rwpos19_75 in19_75 sp19_75 78000.000000
Rwpos19_76 in19_76 sp19_76 78000.000000
Rwpos19_77 in19_77 sp19_77 78000.000000
Rwpos19_78 in19_78 sp19_78 202000.000000
Rwpos19_79 in19_79 sp19_79 78000.000000
Rwpos19_80 in19_80 sp19_80 202000.000000
Rwpos19_81 in19_81 sp19_81 78000.000000
Rwpos19_82 in19_82 sp19_82 78000.000000
Rwpos19_83 in19_83 sp19_83 78000.000000
Rwpos19_84 in19_84 sp19_84 78000.000000
Rwpos20_1 in20_1 sp20_1 202000.000000
Rwpos20_2 in20_2 sp20_2 202000.000000
Rwpos20_3 in20_3 sp20_3 78000.000000
Rwpos20_4 in20_4 sp20_4 202000.000000
Rwpos20_5 in20_5 sp20_5 78000.000000
Rwpos20_6 in20_6 sp20_6 78000.000000
Rwpos20_7 in20_7 sp20_7 202000.000000
Rwpos20_8 in20_8 sp20_8 202000.000000
Rwpos20_9 in20_9 sp20_9 202000.000000
Rwpos20_10 in20_10 sp20_10 78000.000000
Rwpos20_11 in20_11 sp20_11 202000.000000
Rwpos20_12 in20_12 sp20_12 78000.000000
Rwpos20_13 in20_13 sp20_13 78000.000000
Rwpos20_14 in20_14 sp20_14 78000.000000
Rwpos20_15 in20_15 sp20_15 202000.000000
Rwpos20_16 in20_16 sp20_16 78000.000000
Rwpos20_17 in20_17 sp20_17 202000.000000
Rwpos20_18 in20_18 sp20_18 78000.000000
Rwpos20_19 in20_19 sp20_19 202000.000000
Rwpos20_20 in20_20 sp20_20 78000.000000
Rwpos20_21 in20_21 sp20_21 202000.000000
Rwpos20_22 in20_22 sp20_22 78000.000000
Rwpos20_23 in20_23 sp20_23 202000.000000
Rwpos20_24 in20_24 sp20_24 78000.000000
Rwpos20_25 in20_25 sp20_25 202000.000000
Rwpos20_26 in20_26 sp20_26 202000.000000
Rwpos20_27 in20_27 sp20_27 78000.000000
Rwpos20_28 in20_28 sp20_28 78000.000000
Rwpos20_29 in20_29 sp20_29 202000.000000
Rwpos20_30 in20_30 sp20_30 202000.000000
Rwpos20_31 in20_31 sp20_31 202000.000000
Rwpos20_32 in20_32 sp20_32 78000.000000
Rwpos20_33 in20_33 sp20_33 202000.000000
Rwpos20_34 in20_34 sp20_34 202000.000000
Rwpos20_35 in20_35 sp20_35 78000.000000
Rwpos20_36 in20_36 sp20_36 78000.000000
Rwpos20_37 in20_37 sp20_37 202000.000000
Rwpos20_38 in20_38 sp20_38 78000.000000
Rwpos20_39 in20_39 sp20_39 78000.000000
Rwpos20_40 in20_40 sp20_40 202000.000000
Rwpos20_41 in20_41 sp20_41 202000.000000
Rwpos20_42 in20_42 sp20_42 202000.000000
Rwpos20_43 in20_43 sp20_43 202000.000000
Rwpos20_44 in20_44 sp20_44 202000.000000
Rwpos20_45 in20_45 sp20_45 78000.000000
Rwpos20_46 in20_46 sp20_46 202000.000000
Rwpos20_47 in20_47 sp20_47 202000.000000
Rwpos20_48 in20_48 sp20_48 78000.000000
Rwpos20_49 in20_49 sp20_49 202000.000000
Rwpos20_50 in20_50 sp20_50 202000.000000
Rwpos20_51 in20_51 sp20_51 78000.000000
Rwpos20_52 in20_52 sp20_52 202000.000000
Rwpos20_53 in20_53 sp20_53 202000.000000
Rwpos20_54 in20_54 sp20_54 202000.000000
Rwpos20_55 in20_55 sp20_55 202000.000000
Rwpos20_56 in20_56 sp20_56 78000.000000
Rwpos20_57 in20_57 sp20_57 78000.000000
Rwpos20_58 in20_58 sp20_58 202000.000000
Rwpos20_59 in20_59 sp20_59 78000.000000
Rwpos20_60 in20_60 sp20_60 78000.000000
Rwpos20_61 in20_61 sp20_61 78000.000000
Rwpos20_62 in20_62 sp20_62 202000.000000
Rwpos20_63 in20_63 sp20_63 78000.000000
Rwpos20_64 in20_64 sp20_64 202000.000000
Rwpos20_65 in20_65 sp20_65 78000.000000
Rwpos20_66 in20_66 sp20_66 78000.000000
Rwpos20_67 in20_67 sp20_67 78000.000000
Rwpos20_68 in20_68 sp20_68 78000.000000
Rwpos20_69 in20_69 sp20_69 78000.000000
Rwpos20_70 in20_70 sp20_70 78000.000000
Rwpos20_71 in20_71 sp20_71 78000.000000
Rwpos20_72 in20_72 sp20_72 78000.000000
Rwpos20_73 in20_73 sp20_73 78000.000000
Rwpos20_74 in20_74 sp20_74 78000.000000
Rwpos20_75 in20_75 sp20_75 78000.000000
Rwpos20_76 in20_76 sp20_76 202000.000000
Rwpos20_77 in20_77 sp20_77 202000.000000
Rwpos20_78 in20_78 sp20_78 78000.000000
Rwpos20_79 in20_79 sp20_79 78000.000000
Rwpos20_80 in20_80 sp20_80 202000.000000
Rwpos20_81 in20_81 sp20_81 78000.000000
Rwpos20_82 in20_82 sp20_82 78000.000000
Rwpos20_83 in20_83 sp20_83 78000.000000
Rwpos20_84 in20_84 sp20_84 78000.000000
Rwpos21_1 in21_1 sp21_1 202000.000000
Rwpos21_2 in21_2 sp21_2 78000.000000
Rwpos21_3 in21_3 sp21_3 78000.000000
Rwpos21_4 in21_4 sp21_4 78000.000000
Rwpos21_5 in21_5 sp21_5 78000.000000
Rwpos21_6 in21_6 sp21_6 78000.000000
Rwpos21_7 in21_7 sp21_7 78000.000000
Rwpos21_8 in21_8 sp21_8 78000.000000
Rwpos21_9 in21_9 sp21_9 78000.000000
Rwpos21_10 in21_10 sp21_10 78000.000000
Rwpos21_11 in21_11 sp21_11 202000.000000
Rwpos21_12 in21_12 sp21_12 78000.000000
Rwpos21_13 in21_13 sp21_13 78000.000000
Rwpos21_14 in21_14 sp21_14 78000.000000
Rwpos21_15 in21_15 sp21_15 202000.000000
Rwpos21_16 in21_16 sp21_16 202000.000000
Rwpos21_17 in21_17 sp21_17 202000.000000
Rwpos21_18 in21_18 sp21_18 78000.000000
Rwpos21_19 in21_19 sp21_19 202000.000000
Rwpos21_20 in21_20 sp21_20 202000.000000
Rwpos21_21 in21_21 sp21_21 202000.000000
Rwpos21_22 in21_22 sp21_22 202000.000000
Rwpos21_23 in21_23 sp21_23 202000.000000
Rwpos21_24 in21_24 sp21_24 202000.000000
Rwpos21_25 in21_25 sp21_25 202000.000000
Rwpos21_26 in21_26 sp21_26 202000.000000
Rwpos21_27 in21_27 sp21_27 78000.000000
Rwpos21_28 in21_28 sp21_28 202000.000000
Rwpos21_29 in21_29 sp21_29 202000.000000
Rwpos21_30 in21_30 sp21_30 78000.000000
Rwpos21_31 in21_31 sp21_31 202000.000000
Rwpos21_32 in21_32 sp21_32 78000.000000
Rwpos21_33 in21_33 sp21_33 78000.000000
Rwpos21_34 in21_34 sp21_34 202000.000000
Rwpos21_35 in21_35 sp21_35 78000.000000
Rwpos21_36 in21_36 sp21_36 78000.000000
Rwpos21_37 in21_37 sp21_37 202000.000000
Rwpos21_38 in21_38 sp21_38 202000.000000
Rwpos21_39 in21_39 sp21_39 78000.000000
Rwpos21_40 in21_40 sp21_40 202000.000000
Rwpos21_41 in21_41 sp21_41 78000.000000
Rwpos21_42 in21_42 sp21_42 78000.000000
Rwpos21_43 in21_43 sp21_43 78000.000000
Rwpos21_44 in21_44 sp21_44 78000.000000
Rwpos21_45 in21_45 sp21_45 78000.000000
Rwpos21_46 in21_46 sp21_46 202000.000000
Rwpos21_47 in21_47 sp21_47 78000.000000
Rwpos21_48 in21_48 sp21_48 202000.000000
Rwpos21_49 in21_49 sp21_49 78000.000000
Rwpos21_50 in21_50 sp21_50 78000.000000
Rwpos21_51 in21_51 sp21_51 78000.000000
Rwpos21_52 in21_52 sp21_52 78000.000000
Rwpos21_53 in21_53 sp21_53 202000.000000
Rwpos21_54 in21_54 sp21_54 78000.000000
Rwpos21_55 in21_55 sp21_55 78000.000000
Rwpos21_56 in21_56 sp21_56 78000.000000
Rwpos21_57 in21_57 sp21_57 202000.000000
Rwpos21_58 in21_58 sp21_58 202000.000000
Rwpos21_59 in21_59 sp21_59 78000.000000
Rwpos21_60 in21_60 sp21_60 78000.000000
Rwpos21_61 in21_61 sp21_61 78000.000000
Rwpos21_62 in21_62 sp21_62 202000.000000
Rwpos21_63 in21_63 sp21_63 78000.000000
Rwpos21_64 in21_64 sp21_64 78000.000000
Rwpos21_65 in21_65 sp21_65 78000.000000
Rwpos21_66 in21_66 sp21_66 78000.000000
Rwpos21_67 in21_67 sp21_67 202000.000000
Rwpos21_68 in21_68 sp21_68 78000.000000
Rwpos21_69 in21_69 sp21_69 78000.000000
Rwpos21_70 in21_70 sp21_70 202000.000000
Rwpos21_71 in21_71 sp21_71 78000.000000
Rwpos21_72 in21_72 sp21_72 202000.000000
Rwpos21_73 in21_73 sp21_73 202000.000000
Rwpos21_74 in21_74 sp21_74 202000.000000
Rwpos21_75 in21_75 sp21_75 202000.000000
Rwpos21_76 in21_76 sp21_76 78000.000000
Rwpos21_77 in21_77 sp21_77 202000.000000
Rwpos21_78 in21_78 sp21_78 202000.000000
Rwpos21_79 in21_79 sp21_79 78000.000000
Rwpos21_80 in21_80 sp21_80 78000.000000
Rwpos21_81 in21_81 sp21_81 78000.000000
Rwpos21_82 in21_82 sp21_82 78000.000000
Rwpos21_83 in21_83 sp21_83 78000.000000
Rwpos21_84 in21_84 sp21_84 78000.000000
Rwpos22_1 in22_1 sp22_1 202000.000000
Rwpos22_2 in22_2 sp22_2 202000.000000
Rwpos22_3 in22_3 sp22_3 78000.000000
Rwpos22_4 in22_4 sp22_4 78000.000000
Rwpos22_5 in22_5 sp22_5 78000.000000
Rwpos22_6 in22_6 sp22_6 202000.000000
Rwpos22_7 in22_7 sp22_7 78000.000000
Rwpos22_8 in22_8 sp22_8 78000.000000
Rwpos22_9 in22_9 sp22_9 78000.000000
Rwpos22_10 in22_10 sp22_10 202000.000000
Rwpos22_11 in22_11 sp22_11 202000.000000
Rwpos22_12 in22_12 sp22_12 78000.000000
Rwpos22_13 in22_13 sp22_13 78000.000000
Rwpos22_14 in22_14 sp22_14 78000.000000
Rwpos22_15 in22_15 sp22_15 78000.000000
Rwpos22_16 in22_16 sp22_16 78000.000000
Rwpos22_17 in22_17 sp22_17 202000.000000
Rwpos22_18 in22_18 sp22_18 78000.000000
Rwpos22_19 in22_19 sp22_19 202000.000000
Rwpos22_20 in22_20 sp22_20 78000.000000
Rwpos22_21 in22_21 sp22_21 202000.000000
Rwpos22_22 in22_22 sp22_22 78000.000000
Rwpos22_23 in22_23 sp22_23 78000.000000
Rwpos22_24 in22_24 sp22_24 78000.000000
Rwpos22_25 in22_25 sp22_25 202000.000000
Rwpos22_26 in22_26 sp22_26 78000.000000
Rwpos22_27 in22_27 sp22_27 78000.000000
Rwpos22_28 in22_28 sp22_28 78000.000000
Rwpos22_29 in22_29 sp22_29 202000.000000
Rwpos22_30 in22_30 sp22_30 202000.000000
Rwpos22_31 in22_31 sp22_31 202000.000000
Rwpos22_32 in22_32 sp22_32 78000.000000
Rwpos22_33 in22_33 sp22_33 78000.000000
Rwpos22_34 in22_34 sp22_34 78000.000000
Rwpos22_35 in22_35 sp22_35 78000.000000
Rwpos22_36 in22_36 sp22_36 78000.000000
Rwpos22_37 in22_37 sp22_37 202000.000000
Rwpos22_38 in22_38 sp22_38 78000.000000
Rwpos22_39 in22_39 sp22_39 78000.000000
Rwpos22_40 in22_40 sp22_40 202000.000000
Rwpos22_41 in22_41 sp22_41 202000.000000
Rwpos22_42 in22_42 sp22_42 202000.000000
Rwpos22_43 in22_43 sp22_43 202000.000000
Rwpos22_44 in22_44 sp22_44 202000.000000
Rwpos22_45 in22_45 sp22_45 78000.000000
Rwpos22_46 in22_46 sp22_46 78000.000000
Rwpos22_47 in22_47 sp22_47 78000.000000
Rwpos22_48 in22_48 sp22_48 202000.000000
Rwpos22_49 in22_49 sp22_49 78000.000000
Rwpos22_50 in22_50 sp22_50 78000.000000
Rwpos22_51 in22_51 sp22_51 78000.000000
Rwpos22_52 in22_52 sp22_52 78000.000000
Rwpos22_53 in22_53 sp22_53 202000.000000
Rwpos22_54 in22_54 sp22_54 202000.000000
Rwpos22_55 in22_55 sp22_55 202000.000000
Rwpos22_56 in22_56 sp22_56 202000.000000
Rwpos22_57 in22_57 sp22_57 78000.000000
Rwpos22_58 in22_58 sp22_58 202000.000000
Rwpos22_59 in22_59 sp22_59 78000.000000
Rwpos22_60 in22_60 sp22_60 78000.000000
Rwpos22_61 in22_61 sp22_61 202000.000000
Rwpos22_62 in22_62 sp22_62 202000.000000
Rwpos22_63 in22_63 sp22_63 78000.000000
Rwpos22_64 in22_64 sp22_64 202000.000000
Rwpos22_65 in22_65 sp22_65 202000.000000
Rwpos22_66 in22_66 sp22_66 78000.000000
Rwpos22_67 in22_67 sp22_67 78000.000000
Rwpos22_68 in22_68 sp22_68 202000.000000
Rwpos22_69 in22_69 sp22_69 78000.000000
Rwpos22_70 in22_70 sp22_70 78000.000000
Rwpos22_71 in22_71 sp22_71 202000.000000
Rwpos22_72 in22_72 sp22_72 78000.000000
Rwpos22_73 in22_73 sp22_73 202000.000000
Rwpos22_74 in22_74 sp22_74 78000.000000
Rwpos22_75 in22_75 sp22_75 78000.000000
Rwpos22_76 in22_76 sp22_76 78000.000000
Rwpos22_77 in22_77 sp22_77 202000.000000
Rwpos22_78 in22_78 sp22_78 78000.000000
Rwpos22_79 in22_79 sp22_79 78000.000000
Rwpos22_80 in22_80 sp22_80 202000.000000
Rwpos22_81 in22_81 sp22_81 202000.000000
Rwpos22_82 in22_82 sp22_82 78000.000000
Rwpos22_83 in22_83 sp22_83 202000.000000
Rwpos22_84 in22_84 sp22_84 78000.000000
Rwpos23_1 in23_1 sp23_1 78000.000000
Rwpos23_2 in23_2 sp23_2 202000.000000
Rwpos23_3 in23_3 sp23_3 78000.000000
Rwpos23_4 in23_4 sp23_4 78000.000000
Rwpos23_5 in23_5 sp23_5 202000.000000
Rwpos23_6 in23_6 sp23_6 202000.000000
Rwpos23_7 in23_7 sp23_7 78000.000000
Rwpos23_8 in23_8 sp23_8 202000.000000
Rwpos23_9 in23_9 sp23_9 78000.000000
Rwpos23_10 in23_10 sp23_10 202000.000000
Rwpos23_11 in23_11 sp23_11 202000.000000
Rwpos23_12 in23_12 sp23_12 202000.000000
Rwpos23_13 in23_13 sp23_13 202000.000000
Rwpos23_14 in23_14 sp23_14 202000.000000
Rwpos23_15 in23_15 sp23_15 78000.000000
Rwpos23_16 in23_16 sp23_16 202000.000000
Rwpos23_17 in23_17 sp23_17 78000.000000
Rwpos23_18 in23_18 sp23_18 202000.000000
Rwpos23_19 in23_19 sp23_19 202000.000000
Rwpos23_20 in23_20 sp23_20 202000.000000
Rwpos23_21 in23_21 sp23_21 202000.000000
Rwpos23_22 in23_22 sp23_22 202000.000000
Rwpos23_23 in23_23 sp23_23 78000.000000
Rwpos23_24 in23_24 sp23_24 78000.000000
Rwpos23_25 in23_25 sp23_25 78000.000000
Rwpos23_26 in23_26 sp23_26 202000.000000
Rwpos23_27 in23_27 sp23_27 202000.000000
Rwpos23_28 in23_28 sp23_28 202000.000000
Rwpos23_29 in23_29 sp23_29 202000.000000
Rwpos23_30 in23_30 sp23_30 78000.000000
Rwpos23_31 in23_31 sp23_31 202000.000000
Rwpos23_32 in23_32 sp23_32 202000.000000
Rwpos23_33 in23_33 sp23_33 78000.000000
Rwpos23_34 in23_34 sp23_34 78000.000000
Rwpos23_35 in23_35 sp23_35 202000.000000
Rwpos23_36 in23_36 sp23_36 78000.000000
Rwpos23_37 in23_37 sp23_37 78000.000000
Rwpos23_38 in23_38 sp23_38 202000.000000
Rwpos23_39 in23_39 sp23_39 78000.000000
Rwpos23_40 in23_40 sp23_40 202000.000000
Rwpos23_41 in23_41 sp23_41 202000.000000
Rwpos23_42 in23_42 sp23_42 78000.000000
Rwpos23_43 in23_43 sp23_43 202000.000000
Rwpos23_44 in23_44 sp23_44 78000.000000
Rwpos23_45 in23_45 sp23_45 202000.000000
Rwpos23_46 in23_46 sp23_46 202000.000000
Rwpos23_47 in23_47 sp23_47 78000.000000
Rwpos23_48 in23_48 sp23_48 202000.000000
Rwpos23_49 in23_49 sp23_49 78000.000000
Rwpos23_50 in23_50 sp23_50 78000.000000
Rwpos23_51 in23_51 sp23_51 202000.000000
Rwpos23_52 in23_52 sp23_52 78000.000000
Rwpos23_53 in23_53 sp23_53 202000.000000
Rwpos23_54 in23_54 sp23_54 78000.000000
Rwpos23_55 in23_55 sp23_55 202000.000000
Rwpos23_56 in23_56 sp23_56 202000.000000
Rwpos23_57 in23_57 sp23_57 78000.000000
Rwpos23_58 in23_58 sp23_58 202000.000000
Rwpos23_59 in23_59 sp23_59 78000.000000
Rwpos23_60 in23_60 sp23_60 78000.000000
Rwpos23_61 in23_61 sp23_61 202000.000000
Rwpos23_62 in23_62 sp23_62 78000.000000
Rwpos23_63 in23_63 sp23_63 78000.000000
Rwpos23_64 in23_64 sp23_64 202000.000000
Rwpos23_65 in23_65 sp23_65 202000.000000
Rwpos23_66 in23_66 sp23_66 78000.000000
Rwpos23_67 in23_67 sp23_67 202000.000000
Rwpos23_68 in23_68 sp23_68 78000.000000
Rwpos23_69 in23_69 sp23_69 78000.000000
Rwpos23_70 in23_70 sp23_70 78000.000000
Rwpos23_71 in23_71 sp23_71 78000.000000
Rwpos23_72 in23_72 sp23_72 78000.000000
Rwpos23_73 in23_73 sp23_73 78000.000000
Rwpos23_74 in23_74 sp23_74 78000.000000
Rwpos23_75 in23_75 sp23_75 78000.000000
Rwpos23_76 in23_76 sp23_76 78000.000000
Rwpos23_77 in23_77 sp23_77 202000.000000
Rwpos23_78 in23_78 sp23_78 202000.000000
Rwpos23_79 in23_79 sp23_79 78000.000000
Rwpos23_80 in23_80 sp23_80 202000.000000
Rwpos23_81 in23_81 sp23_81 78000.000000
Rwpos23_82 in23_82 sp23_82 78000.000000
Rwpos23_83 in23_83 sp23_83 202000.000000
Rwpos23_84 in23_84 sp23_84 202000.000000
Rwpos24_1 in24_1 sp24_1 202000.000000
Rwpos24_2 in24_2 sp24_2 78000.000000
Rwpos24_3 in24_3 sp24_3 78000.000000
Rwpos24_4 in24_4 sp24_4 202000.000000
Rwpos24_5 in24_5 sp24_5 202000.000000
Rwpos24_6 in24_6 sp24_6 202000.000000
Rwpos24_7 in24_7 sp24_7 78000.000000
Rwpos24_8 in24_8 sp24_8 202000.000000
Rwpos24_9 in24_9 sp24_9 202000.000000
Rwpos24_10 in24_10 sp24_10 78000.000000
Rwpos24_11 in24_11 sp24_11 202000.000000
Rwpos24_12 in24_12 sp24_12 202000.000000
Rwpos24_13 in24_13 sp24_13 78000.000000
Rwpos24_14 in24_14 sp24_14 202000.000000
Rwpos24_15 in24_15 sp24_15 78000.000000
Rwpos24_16 in24_16 sp24_16 202000.000000
Rwpos24_17 in24_17 sp24_17 202000.000000
Rwpos24_18 in24_18 sp24_18 202000.000000
Rwpos24_19 in24_19 sp24_19 202000.000000
Rwpos24_20 in24_20 sp24_20 78000.000000
Rwpos24_21 in24_21 sp24_21 202000.000000
Rwpos24_22 in24_22 sp24_22 202000.000000
Rwpos24_23 in24_23 sp24_23 202000.000000
Rwpos24_24 in24_24 sp24_24 78000.000000
Rwpos24_25 in24_25 sp24_25 202000.000000
Rwpos24_26 in24_26 sp24_26 78000.000000
Rwpos24_27 in24_27 sp24_27 202000.000000
Rwpos24_28 in24_28 sp24_28 202000.000000
Rwpos24_29 in24_29 sp24_29 202000.000000
Rwpos24_30 in24_30 sp24_30 78000.000000
Rwpos24_31 in24_31 sp24_31 202000.000000
Rwpos24_32 in24_32 sp24_32 202000.000000
Rwpos24_33 in24_33 sp24_33 78000.000000
Rwpos24_34 in24_34 sp24_34 202000.000000
Rwpos24_35 in24_35 sp24_35 78000.000000
Rwpos24_36 in24_36 sp24_36 78000.000000
Rwpos24_37 in24_37 sp24_37 78000.000000
Rwpos24_38 in24_38 sp24_38 202000.000000
Rwpos24_39 in24_39 sp24_39 202000.000000
Rwpos24_40 in24_40 sp24_40 202000.000000
Rwpos24_41 in24_41 sp24_41 202000.000000
Rwpos24_42 in24_42 sp24_42 78000.000000
Rwpos24_43 in24_43 sp24_43 78000.000000
Rwpos24_44 in24_44 sp24_44 78000.000000
Rwpos24_45 in24_45 sp24_45 78000.000000
Rwpos24_46 in24_46 sp24_46 202000.000000
Rwpos24_47 in24_47 sp24_47 78000.000000
Rwpos24_48 in24_48 sp24_48 202000.000000
Rwpos24_49 in24_49 sp24_49 202000.000000
Rwpos24_50 in24_50 sp24_50 78000.000000
Rwpos24_51 in24_51 sp24_51 202000.000000
Rwpos24_52 in24_52 sp24_52 78000.000000
Rwpos24_53 in24_53 sp24_53 202000.000000
Rwpos24_54 in24_54 sp24_54 202000.000000
Rwpos24_55 in24_55 sp24_55 78000.000000
Rwpos24_56 in24_56 sp24_56 202000.000000
Rwpos24_57 in24_57 sp24_57 78000.000000
Rwpos24_58 in24_58 sp24_58 202000.000000
Rwpos24_59 in24_59 sp24_59 202000.000000
Rwpos24_60 in24_60 sp24_60 78000.000000
Rwpos24_61 in24_61 sp24_61 202000.000000
Rwpos24_62 in24_62 sp24_62 202000.000000
Rwpos24_63 in24_63 sp24_63 78000.000000
Rwpos24_64 in24_64 sp24_64 202000.000000
Rwpos24_65 in24_65 sp24_65 202000.000000
Rwpos24_66 in24_66 sp24_66 78000.000000
Rwpos24_67 in24_67 sp24_67 202000.000000
Rwpos24_68 in24_68 sp24_68 202000.000000
Rwpos24_69 in24_69 sp24_69 202000.000000
Rwpos24_70 in24_70 sp24_70 78000.000000
Rwpos24_71 in24_71 sp24_71 202000.000000
Rwpos24_72 in24_72 sp24_72 78000.000000
Rwpos24_73 in24_73 sp24_73 202000.000000
Rwpos24_74 in24_74 sp24_74 202000.000000
Rwpos24_75 in24_75 sp24_75 78000.000000
Rwpos24_76 in24_76 sp24_76 78000.000000
Rwpos24_77 in24_77 sp24_77 202000.000000
Rwpos24_78 in24_78 sp24_78 202000.000000
Rwpos24_79 in24_79 sp24_79 202000.000000
Rwpos24_80 in24_80 sp24_80 202000.000000
Rwpos24_81 in24_81 sp24_81 78000.000000
Rwpos24_82 in24_82 sp24_82 78000.000000
Rwpos24_83 in24_83 sp24_83 78000.000000
Rwpos24_84 in24_84 sp24_84 78000.000000
Rwpos25_1 in25_1 sp25_1 78000.000000
Rwpos25_2 in25_2 sp25_2 202000.000000
Rwpos25_3 in25_3 sp25_3 202000.000000
Rwpos25_4 in25_4 sp25_4 202000.000000
Rwpos25_5 in25_5 sp25_5 78000.000000
Rwpos25_6 in25_6 sp25_6 202000.000000
Rwpos25_7 in25_7 sp25_7 78000.000000
Rwpos25_8 in25_8 sp25_8 202000.000000
Rwpos25_9 in25_9 sp25_9 202000.000000
Rwpos25_10 in25_10 sp25_10 78000.000000
Rwpos25_11 in25_11 sp25_11 78000.000000
Rwpos25_12 in25_12 sp25_12 202000.000000
Rwpos25_13 in25_13 sp25_13 78000.000000
Rwpos25_14 in25_14 sp25_14 202000.000000
Rwpos25_15 in25_15 sp25_15 202000.000000
Rwpos25_16 in25_16 sp25_16 78000.000000
Rwpos25_17 in25_17 sp25_17 78000.000000
Rwpos25_18 in25_18 sp25_18 202000.000000
Rwpos25_19 in25_19 sp25_19 78000.000000
Rwpos25_20 in25_20 sp25_20 78000.000000
Rwpos25_21 in25_21 sp25_21 202000.000000
Rwpos25_22 in25_22 sp25_22 78000.000000
Rwpos25_23 in25_23 sp25_23 202000.000000
Rwpos25_24 in25_24 sp25_24 78000.000000
Rwpos25_25 in25_25 sp25_25 78000.000000
Rwpos25_26 in25_26 sp25_26 78000.000000
Rwpos25_27 in25_27 sp25_27 202000.000000
Rwpos25_28 in25_28 sp25_28 78000.000000
Rwpos25_29 in25_29 sp25_29 78000.000000
Rwpos25_30 in25_30 sp25_30 78000.000000
Rwpos25_31 in25_31 sp25_31 202000.000000
Rwpos25_32 in25_32 sp25_32 78000.000000
Rwpos25_33 in25_33 sp25_33 78000.000000
Rwpos25_34 in25_34 sp25_34 78000.000000
Rwpos25_35 in25_35 sp25_35 202000.000000
Rwpos25_36 in25_36 sp25_36 78000.000000
Rwpos25_37 in25_37 sp25_37 78000.000000
Rwpos25_38 in25_38 sp25_38 78000.000000
Rwpos25_39 in25_39 sp25_39 78000.000000
Rwpos25_40 in25_40 sp25_40 78000.000000
Rwpos25_41 in25_41 sp25_41 78000.000000
Rwpos25_42 in25_42 sp25_42 78000.000000
Rwpos25_43 in25_43 sp25_43 78000.000000
Rwpos25_44 in25_44 sp25_44 78000.000000
Rwpos25_45 in25_45 sp25_45 202000.000000
Rwpos25_46 in25_46 sp25_46 202000.000000
Rwpos25_47 in25_47 sp25_47 78000.000000
Rwpos25_48 in25_48 sp25_48 202000.000000
Rwpos25_49 in25_49 sp25_49 78000.000000
Rwpos25_50 in25_50 sp25_50 78000.000000
Rwpos25_51 in25_51 sp25_51 78000.000000
Rwpos25_52 in25_52 sp25_52 78000.000000
Rwpos25_53 in25_53 sp25_53 202000.000000
Rwpos25_54 in25_54 sp25_54 202000.000000
Rwpos25_55 in25_55 sp25_55 78000.000000
Rwpos25_56 in25_56 sp25_56 202000.000000
Rwpos25_57 in25_57 sp25_57 202000.000000
Rwpos25_58 in25_58 sp25_58 78000.000000
Rwpos25_59 in25_59 sp25_59 78000.000000
Rwpos25_60 in25_60 sp25_60 202000.000000
Rwpos25_61 in25_61 sp25_61 202000.000000
Rwpos25_62 in25_62 sp25_62 78000.000000
Rwpos25_63 in25_63 sp25_63 78000.000000
Rwpos25_64 in25_64 sp25_64 202000.000000
Rwpos25_65 in25_65 sp25_65 78000.000000
Rwpos25_66 in25_66 sp25_66 202000.000000
Rwpos25_67 in25_67 sp25_67 78000.000000
Rwpos25_68 in25_68 sp25_68 202000.000000
Rwpos25_69 in25_69 sp25_69 78000.000000
Rwpos25_70 in25_70 sp25_70 78000.000000
Rwpos25_71 in25_71 sp25_71 78000.000000
Rwpos25_72 in25_72 sp25_72 202000.000000
Rwpos25_73 in25_73 sp25_73 202000.000000
Rwpos25_74 in25_74 sp25_74 202000.000000
Rwpos25_75 in25_75 sp25_75 202000.000000
Rwpos25_76 in25_76 sp25_76 202000.000000
Rwpos25_77 in25_77 sp25_77 78000.000000
Rwpos25_78 in25_78 sp25_78 78000.000000
Rwpos25_79 in25_79 sp25_79 78000.000000
Rwpos25_80 in25_80 sp25_80 202000.000000
Rwpos25_81 in25_81 sp25_81 202000.000000
Rwpos25_82 in25_82 sp25_82 202000.000000
Rwpos25_83 in25_83 sp25_83 202000.000000
Rwpos25_84 in25_84 sp25_84 202000.000000
Rwpos26_1 in26_1 sp26_1 78000.000000
Rwpos26_2 in26_2 sp26_2 202000.000000
Rwpos26_3 in26_3 sp26_3 78000.000000
Rwpos26_4 in26_4 sp26_4 78000.000000
Rwpos26_5 in26_5 sp26_5 78000.000000
Rwpos26_6 in26_6 sp26_6 202000.000000
Rwpos26_7 in26_7 sp26_7 202000.000000
Rwpos26_8 in26_8 sp26_8 202000.000000
Rwpos26_9 in26_9 sp26_9 202000.000000
Rwpos26_10 in26_10 sp26_10 202000.000000
Rwpos26_11 in26_11 sp26_11 202000.000000
Rwpos26_12 in26_12 sp26_12 202000.000000
Rwpos26_13 in26_13 sp26_13 202000.000000
Rwpos26_14 in26_14 sp26_14 78000.000000
Rwpos26_15 in26_15 sp26_15 202000.000000
Rwpos26_16 in26_16 sp26_16 202000.000000
Rwpos26_17 in26_17 sp26_17 78000.000000
Rwpos26_18 in26_18 sp26_18 78000.000000
Rwpos26_19 in26_19 sp26_19 202000.000000
Rwpos26_20 in26_20 sp26_20 202000.000000
Rwpos26_21 in26_21 sp26_21 78000.000000
Rwpos26_22 in26_22 sp26_22 78000.000000
Rwpos26_23 in26_23 sp26_23 202000.000000
Rwpos26_24 in26_24 sp26_24 78000.000000
Rwpos26_25 in26_25 sp26_25 78000.000000
Rwpos26_26 in26_26 sp26_26 78000.000000
Rwpos26_27 in26_27 sp26_27 78000.000000
Rwpos26_28 in26_28 sp26_28 78000.000000
Rwpos26_29 in26_29 sp26_29 78000.000000
Rwpos26_30 in26_30 sp26_30 78000.000000
Rwpos26_31 in26_31 sp26_31 202000.000000
Rwpos26_32 in26_32 sp26_32 202000.000000
Rwpos26_33 in26_33 sp26_33 78000.000000
Rwpos26_34 in26_34 sp26_34 202000.000000
Rwpos26_35 in26_35 sp26_35 78000.000000
Rwpos26_36 in26_36 sp26_36 202000.000000
Rwpos26_37 in26_37 sp26_37 202000.000000
Rwpos26_38 in26_38 sp26_38 202000.000000
Rwpos26_39 in26_39 sp26_39 78000.000000
Rwpos26_40 in26_40 sp26_40 202000.000000
Rwpos26_41 in26_41 sp26_41 78000.000000
Rwpos26_42 in26_42 sp26_42 78000.000000
Rwpos26_43 in26_43 sp26_43 202000.000000
Rwpos26_44 in26_44 sp26_44 78000.000000
Rwpos26_45 in26_45 sp26_45 202000.000000
Rwpos26_46 in26_46 sp26_46 78000.000000
Rwpos26_47 in26_47 sp26_47 202000.000000
Rwpos26_48 in26_48 sp26_48 202000.000000
Rwpos26_49 in26_49 sp26_49 202000.000000
Rwpos26_50 in26_50 sp26_50 78000.000000
Rwpos26_51 in26_51 sp26_51 78000.000000
Rwpos26_52 in26_52 sp26_52 202000.000000
Rwpos26_53 in26_53 sp26_53 78000.000000
Rwpos26_54 in26_54 sp26_54 202000.000000
Rwpos26_55 in26_55 sp26_55 202000.000000
Rwpos26_56 in26_56 sp26_56 202000.000000
Rwpos26_57 in26_57 sp26_57 78000.000000
Rwpos26_58 in26_58 sp26_58 202000.000000
Rwpos26_59 in26_59 sp26_59 78000.000000
Rwpos26_60 in26_60 sp26_60 78000.000000
Rwpos26_61 in26_61 sp26_61 78000.000000
Rwpos26_62 in26_62 sp26_62 78000.000000
Rwpos26_63 in26_63 sp26_63 78000.000000
Rwpos26_64 in26_64 sp26_64 78000.000000
Rwpos26_65 in26_65 sp26_65 202000.000000
Rwpos26_66 in26_66 sp26_66 202000.000000
Rwpos26_67 in26_67 sp26_67 78000.000000
Rwpos26_68 in26_68 sp26_68 202000.000000
Rwpos26_69 in26_69 sp26_69 202000.000000
Rwpos26_70 in26_70 sp26_70 202000.000000
Rwpos26_71 in26_71 sp26_71 202000.000000
Rwpos26_72 in26_72 sp26_72 78000.000000
Rwpos26_73 in26_73 sp26_73 202000.000000
Rwpos26_74 in26_74 sp26_74 78000.000000
Rwpos26_75 in26_75 sp26_75 78000.000000
Rwpos26_76 in26_76 sp26_76 202000.000000
Rwpos26_77 in26_77 sp26_77 202000.000000
Rwpos26_78 in26_78 sp26_78 78000.000000
Rwpos26_79 in26_79 sp26_79 202000.000000
Rwpos26_80 in26_80 sp26_80 78000.000000
Rwpos26_81 in26_81 sp26_81 78000.000000
Rwpos26_82 in26_82 sp26_82 78000.000000
Rwpos26_83 in26_83 sp26_83 78000.000000
Rwpos26_84 in26_84 sp26_84 78000.000000
Rwpos27_1 in27_1 sp27_1 78000.000000
Rwpos27_2 in27_2 sp27_2 78000.000000
Rwpos27_3 in27_3 sp27_3 202000.000000
Rwpos27_4 in27_4 sp27_4 78000.000000
Rwpos27_5 in27_5 sp27_5 202000.000000
Rwpos27_6 in27_6 sp27_6 202000.000000
Rwpos27_7 in27_7 sp27_7 78000.000000
Rwpos27_8 in27_8 sp27_8 202000.000000
Rwpos27_9 in27_9 sp27_9 202000.000000
Rwpos27_10 in27_10 sp27_10 202000.000000
Rwpos27_11 in27_11 sp27_11 78000.000000
Rwpos27_12 in27_12 sp27_12 202000.000000
Rwpos27_13 in27_13 sp27_13 202000.000000
Rwpos27_14 in27_14 sp27_14 202000.000000
Rwpos27_15 in27_15 sp27_15 202000.000000
Rwpos27_16 in27_16 sp27_16 78000.000000
Rwpos27_17 in27_17 sp27_17 78000.000000
Rwpos27_18 in27_18 sp27_18 202000.000000
Rwpos27_19 in27_19 sp27_19 78000.000000
Rwpos27_20 in27_20 sp27_20 202000.000000
Rwpos27_21 in27_21 sp27_21 78000.000000
Rwpos27_22 in27_22 sp27_22 78000.000000
Rwpos27_23 in27_23 sp27_23 202000.000000
Rwpos27_24 in27_24 sp27_24 78000.000000
Rwpos27_25 in27_25 sp27_25 78000.000000
Rwpos27_26 in27_26 sp27_26 202000.000000
Rwpos27_27 in27_27 sp27_27 202000.000000
Rwpos27_28 in27_28 sp27_28 78000.000000
Rwpos27_29 in27_29 sp27_29 202000.000000
Rwpos27_30 in27_30 sp27_30 78000.000000
Rwpos27_31 in27_31 sp27_31 202000.000000
Rwpos27_32 in27_32 sp27_32 202000.000000
Rwpos27_33 in27_33 sp27_33 78000.000000
Rwpos27_34 in27_34 sp27_34 202000.000000
Rwpos27_35 in27_35 sp27_35 202000.000000
Rwpos27_36 in27_36 sp27_36 202000.000000
Rwpos27_37 in27_37 sp27_37 78000.000000
Rwpos27_38 in27_38 sp27_38 78000.000000
Rwpos27_39 in27_39 sp27_39 202000.000000
Rwpos27_40 in27_40 sp27_40 78000.000000
Rwpos27_41 in27_41 sp27_41 202000.000000
Rwpos27_42 in27_42 sp27_42 78000.000000
Rwpos27_43 in27_43 sp27_43 202000.000000
Rwpos27_44 in27_44 sp27_44 78000.000000
Rwpos27_45 in27_45 sp27_45 202000.000000
Rwpos27_46 in27_46 sp27_46 202000.000000
Rwpos27_47 in27_47 sp27_47 202000.000000
Rwpos27_48 in27_48 sp27_48 78000.000000
Rwpos27_49 in27_49 sp27_49 78000.000000
Rwpos27_50 in27_50 sp27_50 78000.000000
Rwpos27_51 in27_51 sp27_51 78000.000000
Rwpos27_52 in27_52 sp27_52 78000.000000
Rwpos27_53 in27_53 sp27_53 202000.000000
Rwpos27_54 in27_54 sp27_54 78000.000000
Rwpos27_55 in27_55 sp27_55 78000.000000
Rwpos27_56 in27_56 sp27_56 202000.000000
Rwpos27_57 in27_57 sp27_57 78000.000000
Rwpos27_58 in27_58 sp27_58 78000.000000
Rwpos27_59 in27_59 sp27_59 78000.000000
Rwpos27_60 in27_60 sp27_60 78000.000000
Rwpos27_61 in27_61 sp27_61 78000.000000
Rwpos27_62 in27_62 sp27_62 78000.000000
Rwpos27_63 in27_63 sp27_63 202000.000000
Rwpos27_64 in27_64 sp27_64 78000.000000
Rwpos27_65 in27_65 sp27_65 202000.000000
Rwpos27_66 in27_66 sp27_66 202000.000000
Rwpos27_67 in27_67 sp27_67 202000.000000
Rwpos27_68 in27_68 sp27_68 202000.000000
Rwpos27_69 in27_69 sp27_69 202000.000000
Rwpos27_70 in27_70 sp27_70 202000.000000
Rwpos27_71 in27_71 sp27_71 202000.000000
Rwpos27_72 in27_72 sp27_72 78000.000000
Rwpos27_73 in27_73 sp27_73 78000.000000
Rwpos27_74 in27_74 sp27_74 78000.000000
Rwpos27_75 in27_75 sp27_75 202000.000000
Rwpos27_76 in27_76 sp27_76 202000.000000
Rwpos27_77 in27_77 sp27_77 202000.000000
Rwpos27_78 in27_78 sp27_78 78000.000000
Rwpos27_79 in27_79 sp27_79 202000.000000
Rwpos27_80 in27_80 sp27_80 202000.000000
Rwpos27_81 in27_81 sp27_81 202000.000000
Rwpos27_82 in27_82 sp27_82 202000.000000
Rwpos27_83 in27_83 sp27_83 202000.000000
Rwpos27_84 in27_84 sp27_84 202000.000000
Rwpos28_1 in28_1 sp28_1 78000.000000
Rwpos28_2 in28_2 sp28_2 202000.000000
Rwpos28_3 in28_3 sp28_3 78000.000000
Rwpos28_4 in28_4 sp28_4 78000.000000
Rwpos28_5 in28_5 sp28_5 78000.000000
Rwpos28_6 in28_6 sp28_6 202000.000000
Rwpos28_7 in28_7 sp28_7 202000.000000
Rwpos28_8 in28_8 sp28_8 78000.000000
Rwpos28_9 in28_9 sp28_9 78000.000000
Rwpos28_10 in28_10 sp28_10 202000.000000
Rwpos28_11 in28_11 sp28_11 202000.000000
Rwpos28_12 in28_12 sp28_12 78000.000000
Rwpos28_13 in28_13 sp28_13 202000.000000
Rwpos28_14 in28_14 sp28_14 78000.000000
Rwpos28_15 in28_15 sp28_15 202000.000000
Rwpos28_16 in28_16 sp28_16 78000.000000
Rwpos28_17 in28_17 sp28_17 202000.000000
Rwpos28_18 in28_18 sp28_18 78000.000000
Rwpos28_19 in28_19 sp28_19 202000.000000
Rwpos28_20 in28_20 sp28_20 202000.000000
Rwpos28_21 in28_21 sp28_21 78000.000000
Rwpos28_22 in28_22 sp28_22 202000.000000
Rwpos28_23 in28_23 sp28_23 202000.000000
Rwpos28_24 in28_24 sp28_24 202000.000000
Rwpos28_25 in28_25 sp28_25 78000.000000
Rwpos28_26 in28_26 sp28_26 78000.000000
Rwpos28_27 in28_27 sp28_27 78000.000000
Rwpos28_28 in28_28 sp28_28 78000.000000
Rwpos28_29 in28_29 sp28_29 202000.000000
Rwpos28_30 in28_30 sp28_30 78000.000000
Rwpos28_31 in28_31 sp28_31 78000.000000
Rwpos28_32 in28_32 sp28_32 202000.000000
Rwpos28_33 in28_33 sp28_33 202000.000000
Rwpos28_34 in28_34 sp28_34 78000.000000
Rwpos28_35 in28_35 sp28_35 78000.000000
Rwpos28_36 in28_36 sp28_36 78000.000000
Rwpos28_37 in28_37 sp28_37 78000.000000
Rwpos28_38 in28_38 sp28_38 78000.000000
Rwpos28_39 in28_39 sp28_39 78000.000000
Rwpos28_40 in28_40 sp28_40 202000.000000
Rwpos28_41 in28_41 sp28_41 78000.000000
Rwpos28_42 in28_42 sp28_42 78000.000000
Rwpos28_43 in28_43 sp28_43 78000.000000
Rwpos28_44 in28_44 sp28_44 78000.000000
Rwpos28_45 in28_45 sp28_45 202000.000000
Rwpos28_46 in28_46 sp28_46 78000.000000
Rwpos28_47 in28_47 sp28_47 78000.000000
Rwpos28_48 in28_48 sp28_48 202000.000000
Rwpos28_49 in28_49 sp28_49 78000.000000
Rwpos28_50 in28_50 sp28_50 78000.000000
Rwpos28_51 in28_51 sp28_51 78000.000000
Rwpos28_52 in28_52 sp28_52 78000.000000
Rwpos28_53 in28_53 sp28_53 202000.000000
Rwpos28_54 in28_54 sp28_54 78000.000000
Rwpos28_55 in28_55 sp28_55 202000.000000
Rwpos28_56 in28_56 sp28_56 78000.000000
Rwpos28_57 in28_57 sp28_57 78000.000000
Rwpos28_58 in28_58 sp28_58 202000.000000
Rwpos28_59 in28_59 sp28_59 78000.000000
Rwpos28_60 in28_60 sp28_60 78000.000000
Rwpos28_61 in28_61 sp28_61 78000.000000
Rwpos28_62 in28_62 sp28_62 202000.000000
Rwpos28_63 in28_63 sp28_63 78000.000000
Rwpos28_64 in28_64 sp28_64 202000.000000
Rwpos28_65 in28_65 sp28_65 202000.000000
Rwpos28_66 in28_66 sp28_66 78000.000000
Rwpos28_67 in28_67 sp28_67 78000.000000
Rwpos28_68 in28_68 sp28_68 78000.000000
Rwpos28_69 in28_69 sp28_69 78000.000000
Rwpos28_70 in28_70 sp28_70 202000.000000
Rwpos28_71 in28_71 sp28_71 202000.000000
Rwpos28_72 in28_72 sp28_72 78000.000000
Rwpos28_73 in28_73 sp28_73 78000.000000
Rwpos28_74 in28_74 sp28_74 78000.000000
Rwpos28_75 in28_75 sp28_75 78000.000000
Rwpos28_76 in28_76 sp28_76 78000.000000
Rwpos28_77 in28_77 sp28_77 202000.000000
Rwpos28_78 in28_78 sp28_78 78000.000000
Rwpos28_79 in28_79 sp28_79 78000.000000
Rwpos28_80 in28_80 sp28_80 202000.000000
Rwpos28_81 in28_81 sp28_81 202000.000000
Rwpos28_82 in28_82 sp28_82 78000.000000
Rwpos28_83 in28_83 sp28_83 78000.000000
Rwpos28_84 in28_84 sp28_84 202000.000000
Rwpos29_1 in29_1 sp29_1 202000.000000
Rwpos29_2 in29_2 sp29_2 78000.000000
Rwpos29_3 in29_3 sp29_3 202000.000000
Rwpos29_4 in29_4 sp29_4 202000.000000
Rwpos29_5 in29_5 sp29_5 202000.000000
Rwpos29_6 in29_6 sp29_6 78000.000000
Rwpos29_7 in29_7 sp29_7 202000.000000
Rwpos29_8 in29_8 sp29_8 78000.000000
Rwpos29_9 in29_9 sp29_9 202000.000000
Rwpos29_10 in29_10 sp29_10 202000.000000
Rwpos29_11 in29_11 sp29_11 78000.000000
Rwpos29_12 in29_12 sp29_12 78000.000000
Rwpos29_13 in29_13 sp29_13 78000.000000
Rwpos29_14 in29_14 sp29_14 202000.000000
Rwpos29_15 in29_15 sp29_15 78000.000000
Rwpos29_16 in29_16 sp29_16 78000.000000
Rwpos29_17 in29_17 sp29_17 78000.000000
Rwpos29_18 in29_18 sp29_18 78000.000000
Rwpos29_19 in29_19 sp29_19 78000.000000
Rwpos29_20 in29_20 sp29_20 202000.000000
Rwpos29_21 in29_21 sp29_21 78000.000000
Rwpos29_22 in29_22 sp29_22 78000.000000
Rwpos29_23 in29_23 sp29_23 78000.000000
Rwpos29_24 in29_24 sp29_24 78000.000000
Rwpos29_25 in29_25 sp29_25 202000.000000
Rwpos29_26 in29_26 sp29_26 202000.000000
Rwpos29_27 in29_27 sp29_27 202000.000000
Rwpos29_28 in29_28 sp29_28 202000.000000
Rwpos29_29 in29_29 sp29_29 78000.000000
Rwpos29_30 in29_30 sp29_30 78000.000000
Rwpos29_31 in29_31 sp29_31 78000.000000
Rwpos29_32 in29_32 sp29_32 202000.000000
Rwpos29_33 in29_33 sp29_33 78000.000000
Rwpos29_34 in29_34 sp29_34 202000.000000
Rwpos29_35 in29_35 sp29_35 202000.000000
Rwpos29_36 in29_36 sp29_36 202000.000000
Rwpos29_37 in29_37 sp29_37 202000.000000
Rwpos29_38 in29_38 sp29_38 202000.000000
Rwpos29_39 in29_39 sp29_39 78000.000000
Rwpos29_40 in29_40 sp29_40 202000.000000
Rwpos29_41 in29_41 sp29_41 202000.000000
Rwpos29_42 in29_42 sp29_42 78000.000000
Rwpos29_43 in29_43 sp29_43 202000.000000
Rwpos29_44 in29_44 sp29_44 78000.000000
Rwpos29_45 in29_45 sp29_45 78000.000000
Rwpos29_46 in29_46 sp29_46 202000.000000
Rwpos29_47 in29_47 sp29_47 78000.000000
Rwpos29_48 in29_48 sp29_48 78000.000000
Rwpos29_49 in29_49 sp29_49 202000.000000
Rwpos29_50 in29_50 sp29_50 202000.000000
Rwpos29_51 in29_51 sp29_51 78000.000000
Rwpos29_52 in29_52 sp29_52 202000.000000
Rwpos29_53 in29_53 sp29_53 202000.000000
Rwpos29_54 in29_54 sp29_54 78000.000000
Rwpos29_55 in29_55 sp29_55 78000.000000
Rwpos29_56 in29_56 sp29_56 202000.000000
Rwpos29_57 in29_57 sp29_57 78000.000000
Rwpos29_58 in29_58 sp29_58 202000.000000
Rwpos29_59 in29_59 sp29_59 202000.000000
Rwpos29_60 in29_60 sp29_60 78000.000000
Rwpos29_61 in29_61 sp29_61 78000.000000
Rwpos29_62 in29_62 sp29_62 78000.000000
Rwpos29_63 in29_63 sp29_63 202000.000000
Rwpos29_64 in29_64 sp29_64 78000.000000
Rwpos29_65 in29_65 sp29_65 78000.000000
Rwpos29_66 in29_66 sp29_66 78000.000000
Rwpos29_67 in29_67 sp29_67 202000.000000
Rwpos29_68 in29_68 sp29_68 78000.000000
Rwpos29_69 in29_69 sp29_69 202000.000000
Rwpos29_70 in29_70 sp29_70 78000.000000
Rwpos29_71 in29_71 sp29_71 202000.000000
Rwpos29_72 in29_72 sp29_72 202000.000000
Rwpos29_73 in29_73 sp29_73 78000.000000
Rwpos29_74 in29_74 sp29_74 202000.000000
Rwpos29_75 in29_75 sp29_75 202000.000000
Rwpos29_76 in29_76 sp29_76 202000.000000
Rwpos29_77 in29_77 sp29_77 202000.000000
Rwpos29_78 in29_78 sp29_78 78000.000000
Rwpos29_79 in29_79 sp29_79 202000.000000
Rwpos29_80 in29_80 sp29_80 202000.000000
Rwpos29_81 in29_81 sp29_81 78000.000000
Rwpos29_82 in29_82 sp29_82 202000.000000
Rwpos29_83 in29_83 sp29_83 78000.000000
Rwpos29_84 in29_84 sp29_84 78000.000000
Rwpos30_1 in30_1 sp30_1 78000.000000
Rwpos30_2 in30_2 sp30_2 78000.000000
Rwpos30_3 in30_3 sp30_3 202000.000000
Rwpos30_4 in30_4 sp30_4 202000.000000
Rwpos30_5 in30_5 sp30_5 202000.000000
Rwpos30_6 in30_6 sp30_6 78000.000000
Rwpos30_7 in30_7 sp30_7 202000.000000
Rwpos30_8 in30_8 sp30_8 78000.000000
Rwpos30_9 in30_9 sp30_9 202000.000000
Rwpos30_10 in30_10 sp30_10 78000.000000
Rwpos30_11 in30_11 sp30_11 202000.000000
Rwpos30_12 in30_12 sp30_12 78000.000000
Rwpos30_13 in30_13 sp30_13 78000.000000
Rwpos30_14 in30_14 sp30_14 202000.000000
Rwpos30_15 in30_15 sp30_15 78000.000000
Rwpos30_16 in30_16 sp30_16 78000.000000
Rwpos30_17 in30_17 sp30_17 202000.000000
Rwpos30_18 in30_18 sp30_18 78000.000000
Rwpos30_19 in30_19 sp30_19 78000.000000
Rwpos30_20 in30_20 sp30_20 78000.000000
Rwpos30_21 in30_21 sp30_21 78000.000000
Rwpos30_22 in30_22 sp30_22 78000.000000
Rwpos30_23 in30_23 sp30_23 202000.000000
Rwpos30_24 in30_24 sp30_24 78000.000000
Rwpos30_25 in30_25 sp30_25 78000.000000
Rwpos30_26 in30_26 sp30_26 78000.000000
Rwpos30_27 in30_27 sp30_27 202000.000000
Rwpos30_28 in30_28 sp30_28 78000.000000
Rwpos30_29 in30_29 sp30_29 78000.000000
Rwpos30_30 in30_30 sp30_30 78000.000000
Rwpos30_31 in30_31 sp30_31 202000.000000
Rwpos30_32 in30_32 sp30_32 202000.000000
Rwpos30_33 in30_33 sp30_33 78000.000000
Rwpos30_34 in30_34 sp30_34 202000.000000
Rwpos30_35 in30_35 sp30_35 202000.000000
Rwpos30_36 in30_36 sp30_36 78000.000000
Rwpos30_37 in30_37 sp30_37 202000.000000
Rwpos30_38 in30_38 sp30_38 78000.000000
Rwpos30_39 in30_39 sp30_39 78000.000000
Rwpos30_40 in30_40 sp30_40 78000.000000
Rwpos30_41 in30_41 sp30_41 202000.000000
Rwpos30_42 in30_42 sp30_42 202000.000000
Rwpos30_43 in30_43 sp30_43 202000.000000
Rwpos30_44 in30_44 sp30_44 78000.000000
Rwpos30_45 in30_45 sp30_45 78000.000000
Rwpos30_46 in30_46 sp30_46 202000.000000
Rwpos30_47 in30_47 sp30_47 78000.000000
Rwpos30_48 in30_48 sp30_48 202000.000000
Rwpos30_49 in30_49 sp30_49 78000.000000
Rwpos30_50 in30_50 sp30_50 78000.000000
Rwpos30_51 in30_51 sp30_51 78000.000000
Rwpos30_52 in30_52 sp30_52 202000.000000
Rwpos30_53 in30_53 sp30_53 202000.000000
Rwpos30_54 in30_54 sp30_54 202000.000000
Rwpos30_55 in30_55 sp30_55 78000.000000
Rwpos30_56 in30_56 sp30_56 202000.000000
Rwpos30_57 in30_57 sp30_57 202000.000000
Rwpos30_58 in30_58 sp30_58 202000.000000
Rwpos30_59 in30_59 sp30_59 202000.000000
Rwpos30_60 in30_60 sp30_60 78000.000000
Rwpos30_61 in30_61 sp30_61 78000.000000
Rwpos30_62 in30_62 sp30_62 202000.000000
Rwpos30_63 in30_63 sp30_63 78000.000000
Rwpos30_64 in30_64 sp30_64 202000.000000
Rwpos30_65 in30_65 sp30_65 202000.000000
Rwpos30_66 in30_66 sp30_66 78000.000000
Rwpos30_67 in30_67 sp30_67 78000.000000
Rwpos30_68 in30_68 sp30_68 78000.000000
Rwpos30_69 in30_69 sp30_69 202000.000000
Rwpos30_70 in30_70 sp30_70 202000.000000
Rwpos30_71 in30_71 sp30_71 202000.000000
Rwpos30_72 in30_72 sp30_72 78000.000000
Rwpos30_73 in30_73 sp30_73 202000.000000
Rwpos30_74 in30_74 sp30_74 78000.000000
Rwpos30_75 in30_75 sp30_75 78000.000000
Rwpos30_76 in30_76 sp30_76 202000.000000
Rwpos30_77 in30_77 sp30_77 202000.000000
Rwpos30_78 in30_78 sp30_78 202000.000000
Rwpos30_79 in30_79 sp30_79 202000.000000
Rwpos30_80 in30_80 sp30_80 202000.000000
Rwpos30_81 in30_81 sp30_81 78000.000000
Rwpos30_82 in30_82 sp30_82 78000.000000
Rwpos30_83 in30_83 sp30_83 78000.000000
Rwpos30_84 in30_84 sp30_84 202000.000000
Rwpos31_1 in31_1 sp31_1 78000.000000
Rwpos31_2 in31_2 sp31_2 202000.000000
Rwpos31_3 in31_3 sp31_3 78000.000000
Rwpos31_4 in31_4 sp31_4 78000.000000
Rwpos31_5 in31_5 sp31_5 78000.000000
Rwpos31_6 in31_6 sp31_6 202000.000000
Rwpos31_7 in31_7 sp31_7 202000.000000
Rwpos31_8 in31_8 sp31_8 78000.000000
Rwpos31_9 in31_9 sp31_9 78000.000000
Rwpos31_10 in31_10 sp31_10 78000.000000
Rwpos31_11 in31_11 sp31_11 78000.000000
Rwpos31_12 in31_12 sp31_12 78000.000000
Rwpos31_13 in31_13 sp31_13 78000.000000
Rwpos31_14 in31_14 sp31_14 202000.000000
Rwpos31_15 in31_15 sp31_15 78000.000000
Rwpos31_16 in31_16 sp31_16 202000.000000
Rwpos31_17 in31_17 sp31_17 78000.000000
Rwpos31_18 in31_18 sp31_18 78000.000000
Rwpos31_19 in31_19 sp31_19 202000.000000
Rwpos31_20 in31_20 sp31_20 202000.000000
Rwpos31_21 in31_21 sp31_21 202000.000000
Rwpos31_22 in31_22 sp31_22 78000.000000
Rwpos31_23 in31_23 sp31_23 78000.000000
Rwpos31_24 in31_24 sp31_24 78000.000000
Rwpos31_25 in31_25 sp31_25 78000.000000
Rwpos31_26 in31_26 sp31_26 78000.000000
Rwpos31_27 in31_27 sp31_27 78000.000000
Rwpos31_28 in31_28 sp31_28 202000.000000
Rwpos31_29 in31_29 sp31_29 202000.000000
Rwpos31_30 in31_30 sp31_30 202000.000000
Rwpos31_31 in31_31 sp31_31 78000.000000
Rwpos31_32 in31_32 sp31_32 78000.000000
Rwpos31_33 in31_33 sp31_33 202000.000000
Rwpos31_34 in31_34 sp31_34 78000.000000
Rwpos31_35 in31_35 sp31_35 202000.000000
Rwpos31_36 in31_36 sp31_36 78000.000000
Rwpos31_37 in31_37 sp31_37 202000.000000
Rwpos31_38 in31_38 sp31_38 202000.000000
Rwpos31_39 in31_39 sp31_39 78000.000000
Rwpos31_40 in31_40 sp31_40 202000.000000
Rwpos31_41 in31_41 sp31_41 78000.000000
Rwpos31_42 in31_42 sp31_42 202000.000000
Rwpos31_43 in31_43 sp31_43 202000.000000
Rwpos31_44 in31_44 sp31_44 78000.000000
Rwpos31_45 in31_45 sp31_45 202000.000000
Rwpos31_46 in31_46 sp31_46 202000.000000
Rwpos31_47 in31_47 sp31_47 78000.000000
Rwpos31_48 in31_48 sp31_48 202000.000000
Rwpos31_49 in31_49 sp31_49 78000.000000
Rwpos31_50 in31_50 sp31_50 202000.000000
Rwpos31_51 in31_51 sp31_51 202000.000000
Rwpos31_52 in31_52 sp31_52 202000.000000
Rwpos31_53 in31_53 sp31_53 78000.000000
Rwpos31_54 in31_54 sp31_54 78000.000000
Rwpos31_55 in31_55 sp31_55 202000.000000
Rwpos31_56 in31_56 sp31_56 78000.000000
Rwpos31_57 in31_57 sp31_57 78000.000000
Rwpos31_58 in31_58 sp31_58 78000.000000
Rwpos31_59 in31_59 sp31_59 78000.000000
Rwpos31_60 in31_60 sp31_60 78000.000000
Rwpos31_61 in31_61 sp31_61 78000.000000
Rwpos31_62 in31_62 sp31_62 78000.000000
Rwpos31_63 in31_63 sp31_63 78000.000000
Rwpos31_64 in31_64 sp31_64 202000.000000
Rwpos31_65 in31_65 sp31_65 78000.000000
Rwpos31_66 in31_66 sp31_66 78000.000000
Rwpos31_67 in31_67 sp31_67 202000.000000
Rwpos31_68 in31_68 sp31_68 78000.000000
Rwpos31_69 in31_69 sp31_69 78000.000000
Rwpos31_70 in31_70 sp31_70 202000.000000
Rwpos31_71 in31_71 sp31_71 78000.000000
Rwpos31_72 in31_72 sp31_72 78000.000000
Rwpos31_73 in31_73 sp31_73 78000.000000
Rwpos31_74 in31_74 sp31_74 202000.000000
Rwpos31_75 in31_75 sp31_75 202000.000000
Rwpos31_76 in31_76 sp31_76 78000.000000
Rwpos31_77 in31_77 sp31_77 202000.000000
Rwpos31_78 in31_78 sp31_78 78000.000000
Rwpos31_79 in31_79 sp31_79 78000.000000
Rwpos31_80 in31_80 sp31_80 78000.000000
Rwpos31_81 in31_81 sp31_81 78000.000000
Rwpos31_82 in31_82 sp31_82 78000.000000
Rwpos31_83 in31_83 sp31_83 78000.000000
Rwpos31_84 in31_84 sp31_84 202000.000000
Rwpos32_1 in32_1 sp32_1 202000.000000
Rwpos32_2 in32_2 sp32_2 202000.000000
Rwpos32_3 in32_3 sp32_3 202000.000000
Rwpos32_4 in32_4 sp32_4 78000.000000
Rwpos32_5 in32_5 sp32_5 78000.000000
Rwpos32_6 in32_6 sp32_6 78000.000000
Rwpos32_7 in32_7 sp32_7 202000.000000
Rwpos32_8 in32_8 sp32_8 78000.000000
Rwpos32_9 in32_9 sp32_9 78000.000000
Rwpos32_10 in32_10 sp32_10 202000.000000
Rwpos32_11 in32_11 sp32_11 78000.000000
Rwpos32_12 in32_12 sp32_12 202000.000000
Rwpos32_13 in32_13 sp32_13 78000.000000
Rwpos32_14 in32_14 sp32_14 78000.000000
Rwpos32_15 in32_15 sp32_15 78000.000000
Rwpos32_16 in32_16 sp32_16 78000.000000
Rwpos32_17 in32_17 sp32_17 78000.000000
Rwpos32_18 in32_18 sp32_18 202000.000000
Rwpos32_19 in32_19 sp32_19 78000.000000
Rwpos32_20 in32_20 sp32_20 202000.000000
Rwpos32_21 in32_21 sp32_21 78000.000000
Rwpos32_22 in32_22 sp32_22 78000.000000
Rwpos32_23 in32_23 sp32_23 78000.000000
Rwpos32_24 in32_24 sp32_24 202000.000000
Rwpos32_25 in32_25 sp32_25 202000.000000
Rwpos32_26 in32_26 sp32_26 78000.000000
Rwpos32_27 in32_27 sp32_27 78000.000000
Rwpos32_28 in32_28 sp32_28 202000.000000
Rwpos32_29 in32_29 sp32_29 202000.000000
Rwpos32_30 in32_30 sp32_30 78000.000000
Rwpos32_31 in32_31 sp32_31 78000.000000
Rwpos32_32 in32_32 sp32_32 78000.000000
Rwpos32_33 in32_33 sp32_33 202000.000000
Rwpos32_34 in32_34 sp32_34 202000.000000
Rwpos32_35 in32_35 sp32_35 78000.000000
Rwpos32_36 in32_36 sp32_36 202000.000000
Rwpos32_37 in32_37 sp32_37 78000.000000
Rwpos32_38 in32_38 sp32_38 202000.000000
Rwpos32_39 in32_39 sp32_39 78000.000000
Rwpos32_40 in32_40 sp32_40 78000.000000
Rwpos32_41 in32_41 sp32_41 202000.000000
Rwpos32_42 in32_42 sp32_42 78000.000000
Rwpos32_43 in32_43 sp32_43 78000.000000
Rwpos32_44 in32_44 sp32_44 202000.000000
Rwpos32_45 in32_45 sp32_45 202000.000000
Rwpos32_46 in32_46 sp32_46 78000.000000
Rwpos32_47 in32_47 sp32_47 202000.000000
Rwpos32_48 in32_48 sp32_48 202000.000000
Rwpos32_49 in32_49 sp32_49 202000.000000
Rwpos32_50 in32_50 sp32_50 202000.000000
Rwpos32_51 in32_51 sp32_51 202000.000000
Rwpos32_52 in32_52 sp32_52 202000.000000
Rwpos32_53 in32_53 sp32_53 202000.000000
Rwpos32_54 in32_54 sp32_54 78000.000000
Rwpos32_55 in32_55 sp32_55 202000.000000
Rwpos32_56 in32_56 sp32_56 202000.000000
Rwpos32_57 in32_57 sp32_57 202000.000000
Rwpos32_58 in32_58 sp32_58 78000.000000
Rwpos32_59 in32_59 sp32_59 78000.000000
Rwpos32_60 in32_60 sp32_60 202000.000000
Rwpos32_61 in32_61 sp32_61 202000.000000
Rwpos32_62 in32_62 sp32_62 78000.000000
Rwpos32_63 in32_63 sp32_63 78000.000000
Rwpos32_64 in32_64 sp32_64 202000.000000
Rwpos32_65 in32_65 sp32_65 202000.000000
Rwpos32_66 in32_66 sp32_66 202000.000000
Rwpos32_67 in32_67 sp32_67 78000.000000
Rwpos32_68 in32_68 sp32_68 202000.000000
Rwpos32_69 in32_69 sp32_69 78000.000000
Rwpos32_70 in32_70 sp32_70 78000.000000
Rwpos32_71 in32_71 sp32_71 202000.000000
Rwpos32_72 in32_72 sp32_72 202000.000000
Rwpos32_73 in32_73 sp32_73 202000.000000
Rwpos32_74 in32_74 sp32_74 202000.000000
Rwpos32_75 in32_75 sp32_75 202000.000000
Rwpos32_76 in32_76 sp32_76 202000.000000
Rwpos32_77 in32_77 sp32_77 78000.000000
Rwpos32_78 in32_78 sp32_78 78000.000000
Rwpos32_79 in32_79 sp32_79 78000.000000
Rwpos32_80 in32_80 sp32_80 78000.000000
Rwpos32_81 in32_81 sp32_81 78000.000000
Rwpos32_82 in32_82 sp32_82 202000.000000
Rwpos32_83 in32_83 sp32_83 78000.000000
Rwpos32_84 in32_84 sp32_84 78000.000000
Rwpos33_1 in33_1 sp33_1 202000.000000
Rwpos33_2 in33_2 sp33_2 202000.000000
Rwpos33_3 in33_3 sp33_3 78000.000000
Rwpos33_4 in33_4 sp33_4 78000.000000
Rwpos33_5 in33_5 sp33_5 78000.000000
Rwpos33_6 in33_6 sp33_6 78000.000000
Rwpos33_7 in33_7 sp33_7 202000.000000
Rwpos33_8 in33_8 sp33_8 78000.000000
Rwpos33_9 in33_9 sp33_9 202000.000000
Rwpos33_10 in33_10 sp33_10 202000.000000
Rwpos33_11 in33_11 sp33_11 202000.000000
Rwpos33_12 in33_12 sp33_12 78000.000000
Rwpos33_13 in33_13 sp33_13 78000.000000
Rwpos33_14 in33_14 sp33_14 202000.000000
Rwpos33_15 in33_15 sp33_15 78000.000000
Rwpos33_16 in33_16 sp33_16 202000.000000
Rwpos33_17 in33_17 sp33_17 78000.000000
Rwpos33_18 in33_18 sp33_18 78000.000000
Rwpos33_19 in33_19 sp33_19 78000.000000
Rwpos33_20 in33_20 sp33_20 78000.000000
Rwpos33_21 in33_21 sp33_21 78000.000000
Rwpos33_22 in33_22 sp33_22 78000.000000
Rwpos33_23 in33_23 sp33_23 78000.000000
Rwpos33_24 in33_24 sp33_24 78000.000000
Rwpos33_25 in33_25 sp33_25 78000.000000
Rwpos33_26 in33_26 sp33_26 202000.000000
Rwpos33_27 in33_27 sp33_27 202000.000000
Rwpos33_28 in33_28 sp33_28 78000.000000
Rwpos33_29 in33_29 sp33_29 202000.000000
Rwpos33_30 in33_30 sp33_30 78000.000000
Rwpos33_31 in33_31 sp33_31 202000.000000
Rwpos33_32 in33_32 sp33_32 202000.000000
Rwpos33_33 in33_33 sp33_33 78000.000000
Rwpos33_34 in33_34 sp33_34 202000.000000
Rwpos33_35 in33_35 sp33_35 202000.000000
Rwpos33_36 in33_36 sp33_36 78000.000000
Rwpos33_37 in33_37 sp33_37 202000.000000
Rwpos33_38 in33_38 sp33_38 78000.000000
Rwpos33_39 in33_39 sp33_39 78000.000000
Rwpos33_40 in33_40 sp33_40 78000.000000
Rwpos33_41 in33_41 sp33_41 78000.000000
Rwpos33_42 in33_42 sp33_42 202000.000000
Rwpos33_43 in33_43 sp33_43 78000.000000
Rwpos33_44 in33_44 sp33_44 78000.000000
Rwpos33_45 in33_45 sp33_45 78000.000000
Rwpos33_46 in33_46 sp33_46 202000.000000
Rwpos33_47 in33_47 sp33_47 78000.000000
Rwpos33_48 in33_48 sp33_48 78000.000000
Rwpos33_49 in33_49 sp33_49 202000.000000
Rwpos33_50 in33_50 sp33_50 202000.000000
Rwpos33_51 in33_51 sp33_51 202000.000000
Rwpos33_52 in33_52 sp33_52 202000.000000
Rwpos33_53 in33_53 sp33_53 78000.000000
Rwpos33_54 in33_54 sp33_54 78000.000000
Rwpos33_55 in33_55 sp33_55 202000.000000
Rwpos33_56 in33_56 sp33_56 202000.000000
Rwpos33_57 in33_57 sp33_57 78000.000000
Rwpos33_58 in33_58 sp33_58 78000.000000
Rwpos33_59 in33_59 sp33_59 202000.000000
Rwpos33_60 in33_60 sp33_60 78000.000000
Rwpos33_61 in33_61 sp33_61 78000.000000
Rwpos33_62 in33_62 sp33_62 78000.000000
Rwpos33_63 in33_63 sp33_63 78000.000000
Rwpos33_64 in33_64 sp33_64 78000.000000
Rwpos33_65 in33_65 sp33_65 202000.000000
Rwpos33_66 in33_66 sp33_66 78000.000000
Rwpos33_67 in33_67 sp33_67 78000.000000
Rwpos33_68 in33_68 sp33_68 78000.000000
Rwpos33_69 in33_69 sp33_69 202000.000000
Rwpos33_70 in33_70 sp33_70 78000.000000
Rwpos33_71 in33_71 sp33_71 78000.000000
Rwpos33_72 in33_72 sp33_72 202000.000000
Rwpos33_73 in33_73 sp33_73 202000.000000
Rwpos33_74 in33_74 sp33_74 202000.000000
Rwpos33_75 in33_75 sp33_75 78000.000000
Rwpos33_76 in33_76 sp33_76 202000.000000
Rwpos33_77 in33_77 sp33_77 78000.000000
Rwpos33_78 in33_78 sp33_78 202000.000000
Rwpos33_79 in33_79 sp33_79 78000.000000
Rwpos33_80 in33_80 sp33_80 202000.000000
Rwpos33_81 in33_81 sp33_81 78000.000000
Rwpos33_82 in33_82 sp33_82 202000.000000
Rwpos33_83 in33_83 sp33_83 78000.000000
Rwpos33_84 in33_84 sp33_84 78000.000000
Rwpos34_1 in34_1 sp34_1 78000.000000
Rwpos34_2 in34_2 sp34_2 202000.000000
Rwpos34_3 in34_3 sp34_3 202000.000000
Rwpos34_4 in34_4 sp34_4 202000.000000
Rwpos34_5 in34_5 sp34_5 202000.000000
Rwpos34_6 in34_6 sp34_6 78000.000000
Rwpos34_7 in34_7 sp34_7 202000.000000
Rwpos34_8 in34_8 sp34_8 202000.000000
Rwpos34_9 in34_9 sp34_9 202000.000000
Rwpos34_10 in34_10 sp34_10 78000.000000
Rwpos34_11 in34_11 sp34_11 78000.000000
Rwpos34_12 in34_12 sp34_12 78000.000000
Rwpos34_13 in34_13 sp34_13 78000.000000
Rwpos34_14 in34_14 sp34_14 202000.000000
Rwpos34_15 in34_15 sp34_15 78000.000000
Rwpos34_16 in34_16 sp34_16 78000.000000
Rwpos34_17 in34_17 sp34_17 202000.000000
Rwpos34_18 in34_18 sp34_18 78000.000000
Rwpos34_19 in34_19 sp34_19 78000.000000
Rwpos34_20 in34_20 sp34_20 78000.000000
Rwpos34_21 in34_21 sp34_21 78000.000000
Rwpos34_22 in34_22 sp34_22 78000.000000
Rwpos34_23 in34_23 sp34_23 202000.000000
Rwpos34_24 in34_24 sp34_24 78000.000000
Rwpos34_25 in34_25 sp34_25 78000.000000
Rwpos34_26 in34_26 sp34_26 78000.000000
Rwpos34_27 in34_27 sp34_27 202000.000000
Rwpos34_28 in34_28 sp34_28 78000.000000
Rwpos34_29 in34_29 sp34_29 202000.000000
Rwpos34_30 in34_30 sp34_30 78000.000000
Rwpos34_31 in34_31 sp34_31 202000.000000
Rwpos34_32 in34_32 sp34_32 78000.000000
Rwpos34_33 in34_33 sp34_33 78000.000000
Rwpos34_34 in34_34 sp34_34 78000.000000
Rwpos34_35 in34_35 sp34_35 202000.000000
Rwpos34_36 in34_36 sp34_36 78000.000000
Rwpos34_37 in34_37 sp34_37 202000.000000
Rwpos34_38 in34_38 sp34_38 78000.000000
Rwpos34_39 in34_39 sp34_39 78000.000000
Rwpos34_40 in34_40 sp34_40 78000.000000
Rwpos34_41 in34_41 sp34_41 202000.000000
Rwpos34_42 in34_42 sp34_42 202000.000000
Rwpos34_43 in34_43 sp34_43 202000.000000
Rwpos34_44 in34_44 sp34_44 78000.000000
Rwpos34_45 in34_45 sp34_45 78000.000000
Rwpos34_46 in34_46 sp34_46 202000.000000
Rwpos34_47 in34_47 sp34_47 78000.000000
Rwpos34_48 in34_48 sp34_48 202000.000000
Rwpos34_49 in34_49 sp34_49 78000.000000
Rwpos34_50 in34_50 sp34_50 202000.000000
Rwpos34_51 in34_51 sp34_51 78000.000000
Rwpos34_52 in34_52 sp34_52 202000.000000
Rwpos34_53 in34_53 sp34_53 202000.000000
Rwpos34_54 in34_54 sp34_54 78000.000000
Rwpos34_55 in34_55 sp34_55 202000.000000
Rwpos34_56 in34_56 sp34_56 78000.000000
Rwpos34_57 in34_57 sp34_57 78000.000000
Rwpos34_58 in34_58 sp34_58 202000.000000
Rwpos34_59 in34_59 sp34_59 78000.000000
Rwpos34_60 in34_60 sp34_60 202000.000000
Rwpos34_61 in34_61 sp34_61 202000.000000
Rwpos34_62 in34_62 sp34_62 202000.000000
Rwpos34_63 in34_63 sp34_63 78000.000000
Rwpos34_64 in34_64 sp34_64 78000.000000
Rwpos34_65 in34_65 sp34_65 78000.000000
Rwpos34_66 in34_66 sp34_66 202000.000000
Rwpos34_67 in34_67 sp34_67 78000.000000
Rwpos34_68 in34_68 sp34_68 78000.000000
Rwpos34_69 in34_69 sp34_69 78000.000000
Rwpos34_70 in34_70 sp34_70 202000.000000
Rwpos34_71 in34_71 sp34_71 78000.000000
Rwpos34_72 in34_72 sp34_72 78000.000000
Rwpos34_73 in34_73 sp34_73 202000.000000
Rwpos34_74 in34_74 sp34_74 202000.000000
Rwpos34_75 in34_75 sp34_75 78000.000000
Rwpos34_76 in34_76 sp34_76 202000.000000
Rwpos34_77 in34_77 sp34_77 78000.000000
Rwpos34_78 in34_78 sp34_78 78000.000000
Rwpos34_79 in34_79 sp34_79 78000.000000
Rwpos34_80 in34_80 sp34_80 202000.000000
Rwpos34_81 in34_81 sp34_81 202000.000000
Rwpos34_82 in34_82 sp34_82 78000.000000
Rwpos34_83 in34_83 sp34_83 202000.000000
Rwpos34_84 in34_84 sp34_84 202000.000000
Rwpos35_1 in35_1 sp35_1 78000.000000
Rwpos35_2 in35_2 sp35_2 78000.000000
Rwpos35_3 in35_3 sp35_3 78000.000000
Rwpos35_4 in35_4 sp35_4 202000.000000
Rwpos35_5 in35_5 sp35_5 78000.000000
Rwpos35_6 in35_6 sp35_6 78000.000000
Rwpos35_7 in35_7 sp35_7 78000.000000
Rwpos35_8 in35_8 sp35_8 202000.000000
Rwpos35_9 in35_9 sp35_9 78000.000000
Rwpos35_10 in35_10 sp35_10 78000.000000
Rwpos35_11 in35_11 sp35_11 78000.000000
Rwpos35_12 in35_12 sp35_12 202000.000000
Rwpos35_13 in35_13 sp35_13 202000.000000
Rwpos35_14 in35_14 sp35_14 78000.000000
Rwpos35_15 in35_15 sp35_15 78000.000000
Rwpos35_16 in35_16 sp35_16 78000.000000
Rwpos35_17 in35_17 sp35_17 78000.000000
Rwpos35_18 in35_18 sp35_18 202000.000000
Rwpos35_19 in35_19 sp35_19 78000.000000
Rwpos35_20 in35_20 sp35_20 78000.000000
Rwpos35_21 in35_21 sp35_21 78000.000000
Rwpos35_22 in35_22 sp35_22 78000.000000
Rwpos35_23 in35_23 sp35_23 202000.000000
Rwpos35_24 in35_24 sp35_24 78000.000000
Rwpos35_25 in35_25 sp35_25 202000.000000
Rwpos35_26 in35_26 sp35_26 202000.000000
Rwpos35_27 in35_27 sp35_27 202000.000000
Rwpos35_28 in35_28 sp35_28 78000.000000
Rwpos35_29 in35_29 sp35_29 78000.000000
Rwpos35_30 in35_30 sp35_30 202000.000000
Rwpos35_31 in35_31 sp35_31 202000.000000
Rwpos35_32 in35_32 sp35_32 78000.000000
Rwpos35_33 in35_33 sp35_33 78000.000000
Rwpos35_34 in35_34 sp35_34 202000.000000
Rwpos35_35 in35_35 sp35_35 202000.000000
Rwpos35_36 in35_36 sp35_36 202000.000000
Rwpos35_37 in35_37 sp35_37 78000.000000
Rwpos35_38 in35_38 sp35_38 78000.000000
Rwpos35_39 in35_39 sp35_39 202000.000000
Rwpos35_40 in35_40 sp35_40 78000.000000
Rwpos35_41 in35_41 sp35_41 78000.000000
Rwpos35_42 in35_42 sp35_42 78000.000000
Rwpos35_43 in35_43 sp35_43 78000.000000
Rwpos35_44 in35_44 sp35_44 78000.000000
Rwpos35_45 in35_45 sp35_45 78000.000000
Rwpos35_46 in35_46 sp35_46 202000.000000
Rwpos35_47 in35_47 sp35_47 78000.000000
Rwpos35_48 in35_48 sp35_48 202000.000000
Rwpos35_49 in35_49 sp35_49 78000.000000
Rwpos35_50 in35_50 sp35_50 78000.000000
Rwpos35_51 in35_51 sp35_51 78000.000000
Rwpos35_52 in35_52 sp35_52 78000.000000
Rwpos35_53 in35_53 sp35_53 202000.000000
Rwpos35_54 in35_54 sp35_54 202000.000000
Rwpos35_55 in35_55 sp35_55 202000.000000
Rwpos35_56 in35_56 sp35_56 202000.000000
Rwpos35_57 in35_57 sp35_57 78000.000000
Rwpos35_58 in35_58 sp35_58 78000.000000
Rwpos35_59 in35_59 sp35_59 202000.000000
Rwpos35_60 in35_60 sp35_60 202000.000000
Rwpos35_61 in35_61 sp35_61 202000.000000
Rwpos35_62 in35_62 sp35_62 78000.000000
Rwpos35_63 in35_63 sp35_63 202000.000000
Rwpos35_64 in35_64 sp35_64 202000.000000
Rwpos35_65 in35_65 sp35_65 202000.000000
Rwpos35_66 in35_66 sp35_66 78000.000000
Rwpos35_67 in35_67 sp35_67 202000.000000
Rwpos35_68 in35_68 sp35_68 202000.000000
Rwpos35_69 in35_69 sp35_69 202000.000000
Rwpos35_70 in35_70 sp35_70 202000.000000
Rwpos35_71 in35_71 sp35_71 202000.000000
Rwpos35_72 in35_72 sp35_72 78000.000000
Rwpos35_73 in35_73 sp35_73 202000.000000
Rwpos35_74 in35_74 sp35_74 202000.000000
Rwpos35_75 in35_75 sp35_75 78000.000000
Rwpos35_76 in35_76 sp35_76 202000.000000
Rwpos35_77 in35_77 sp35_77 202000.000000
Rwpos35_78 in35_78 sp35_78 78000.000000
Rwpos35_79 in35_79 sp35_79 202000.000000
Rwpos35_80 in35_80 sp35_80 202000.000000
Rwpos35_81 in35_81 sp35_81 202000.000000
Rwpos35_82 in35_82 sp35_82 202000.000000
Rwpos35_83 in35_83 sp35_83 202000.000000
Rwpos35_84 in35_84 sp35_84 202000.000000
Rwpos36_1 in36_1 sp36_1 78000.000000
Rwpos36_2 in36_2 sp36_2 78000.000000
Rwpos36_3 in36_3 sp36_3 78000.000000
Rwpos36_4 in36_4 sp36_4 202000.000000
Rwpos36_5 in36_5 sp36_5 202000.000000
Rwpos36_6 in36_6 sp36_6 202000.000000
Rwpos36_7 in36_7 sp36_7 78000.000000
Rwpos36_8 in36_8 sp36_8 78000.000000
Rwpos36_9 in36_9 sp36_9 202000.000000
Rwpos36_10 in36_10 sp36_10 78000.000000
Rwpos36_11 in36_11 sp36_11 202000.000000
Rwpos36_12 in36_12 sp36_12 202000.000000
Rwpos36_13 in36_13 sp36_13 202000.000000
Rwpos36_14 in36_14 sp36_14 202000.000000
Rwpos36_15 in36_15 sp36_15 202000.000000
Rwpos36_16 in36_16 sp36_16 202000.000000
Rwpos36_17 in36_17 sp36_17 202000.000000
Rwpos36_18 in36_18 sp36_18 202000.000000
Rwpos36_19 in36_19 sp36_19 202000.000000
Rwpos36_20 in36_20 sp36_20 78000.000000
Rwpos36_21 in36_21 sp36_21 202000.000000
Rwpos36_22 in36_22 sp36_22 202000.000000
Rwpos36_23 in36_23 sp36_23 78000.000000
Rwpos36_24 in36_24 sp36_24 78000.000000
Rwpos36_25 in36_25 sp36_25 78000.000000
Rwpos36_26 in36_26 sp36_26 78000.000000
Rwpos36_27 in36_27 sp36_27 202000.000000
Rwpos36_28 in36_28 sp36_28 78000.000000
Rwpos36_29 in36_29 sp36_29 78000.000000
Rwpos36_30 in36_30 sp36_30 202000.000000
Rwpos36_31 in36_31 sp36_31 202000.000000
Rwpos36_32 in36_32 sp36_32 202000.000000
Rwpos36_33 in36_33 sp36_33 78000.000000
Rwpos36_34 in36_34 sp36_34 202000.000000
Rwpos36_35 in36_35 sp36_35 78000.000000
Rwpos36_36 in36_36 sp36_36 78000.000000
Rwpos36_37 in36_37 sp36_37 78000.000000
Rwpos36_38 in36_38 sp36_38 202000.000000
Rwpos36_39 in36_39 sp36_39 202000.000000
Rwpos36_40 in36_40 sp36_40 202000.000000
Rwpos36_41 in36_41 sp36_41 202000.000000
Rwpos36_42 in36_42 sp36_42 78000.000000
Rwpos36_43 in36_43 sp36_43 78000.000000
Rwpos36_44 in36_44 sp36_44 78000.000000
Rwpos36_45 in36_45 sp36_45 202000.000000
Rwpos36_46 in36_46 sp36_46 78000.000000
Rwpos36_47 in36_47 sp36_47 78000.000000
Rwpos36_48 in36_48 sp36_48 78000.000000
Rwpos36_49 in36_49 sp36_49 78000.000000
Rwpos36_50 in36_50 sp36_50 78000.000000
Rwpos36_51 in36_51 sp36_51 78000.000000
Rwpos36_52 in36_52 sp36_52 78000.000000
Rwpos36_53 in36_53 sp36_53 78000.000000
Rwpos36_54 in36_54 sp36_54 202000.000000
Rwpos36_55 in36_55 sp36_55 202000.000000
Rwpos36_56 in36_56 sp36_56 78000.000000
Rwpos36_57 in36_57 sp36_57 202000.000000
Rwpos36_58 in36_58 sp36_58 202000.000000
Rwpos36_59 in36_59 sp36_59 202000.000000
Rwpos36_60 in36_60 sp36_60 78000.000000
Rwpos36_61 in36_61 sp36_61 78000.000000
Rwpos36_62 in36_62 sp36_62 78000.000000
Rwpos36_63 in36_63 sp36_63 78000.000000
Rwpos36_64 in36_64 sp36_64 202000.000000
Rwpos36_65 in36_65 sp36_65 78000.000000
Rwpos36_66 in36_66 sp36_66 78000.000000
Rwpos36_67 in36_67 sp36_67 202000.000000
Rwpos36_68 in36_68 sp36_68 202000.000000
Rwpos36_69 in36_69 sp36_69 78000.000000
Rwpos36_70 in36_70 sp36_70 78000.000000
Rwpos36_71 in36_71 sp36_71 78000.000000
Rwpos36_72 in36_72 sp36_72 78000.000000
Rwpos36_73 in36_73 sp36_73 202000.000000
Rwpos36_74 in36_74 sp36_74 202000.000000
Rwpos36_75 in36_75 sp36_75 202000.000000
Rwpos36_76 in36_76 sp36_76 78000.000000
Rwpos36_77 in36_77 sp36_77 202000.000000
Rwpos36_78 in36_78 sp36_78 78000.000000
Rwpos36_79 in36_79 sp36_79 78000.000000
Rwpos36_80 in36_80 sp36_80 202000.000000
Rwpos36_81 in36_81 sp36_81 78000.000000
Rwpos36_82 in36_82 sp36_82 78000.000000
Rwpos36_83 in36_83 sp36_83 202000.000000
Rwpos36_84 in36_84 sp36_84 202000.000000
Rwpos37_1 in37_1 sp37_1 78000.000000
Rwpos37_2 in37_2 sp37_2 202000.000000
Rwpos37_3 in37_3 sp37_3 78000.000000
Rwpos37_4 in37_4 sp37_4 202000.000000
Rwpos37_5 in37_5 sp37_5 78000.000000
Rwpos37_6 in37_6 sp37_6 78000.000000
Rwpos37_7 in37_7 sp37_7 202000.000000
Rwpos37_8 in37_8 sp37_8 202000.000000
Rwpos37_9 in37_9 sp37_9 78000.000000
Rwpos37_10 in37_10 sp37_10 78000.000000
Rwpos37_11 in37_11 sp37_11 202000.000000
Rwpos37_12 in37_12 sp37_12 78000.000000
Rwpos37_13 in37_13 sp37_13 78000.000000
Rwpos37_14 in37_14 sp37_14 78000.000000
Rwpos37_15 in37_15 sp37_15 78000.000000
Rwpos37_16 in37_16 sp37_16 78000.000000
Rwpos37_17 in37_17 sp37_17 202000.000000
Rwpos37_18 in37_18 sp37_18 78000.000000
Rwpos37_19 in37_19 sp37_19 78000.000000
Rwpos37_20 in37_20 sp37_20 78000.000000
Rwpos37_21 in37_21 sp37_21 78000.000000
Rwpos37_22 in37_22 sp37_22 78000.000000
Rwpos37_23 in37_23 sp37_23 202000.000000
Rwpos37_24 in37_24 sp37_24 78000.000000
Rwpos37_25 in37_25 sp37_25 202000.000000
Rwpos37_26 in37_26 sp37_26 202000.000000
Rwpos37_27 in37_27 sp37_27 78000.000000
Rwpos37_28 in37_28 sp37_28 78000.000000
Rwpos37_29 in37_29 sp37_29 78000.000000
Rwpos37_30 in37_30 sp37_30 78000.000000
Rwpos37_31 in37_31 sp37_31 78000.000000
Rwpos37_32 in37_32 sp37_32 202000.000000
Rwpos37_33 in37_33 sp37_33 202000.000000
Rwpos37_34 in37_34 sp37_34 78000.000000
Rwpos37_35 in37_35 sp37_35 78000.000000
Rwpos37_36 in37_36 sp37_36 78000.000000
Rwpos37_37 in37_37 sp37_37 202000.000000
Rwpos37_38 in37_38 sp37_38 78000.000000
Rwpos37_39 in37_39 sp37_39 78000.000000
Rwpos37_40 in37_40 sp37_40 78000.000000
Rwpos37_41 in37_41 sp37_41 202000.000000
Rwpos37_42 in37_42 sp37_42 202000.000000
Rwpos37_43 in37_43 sp37_43 202000.000000
Rwpos37_44 in37_44 sp37_44 202000.000000
Rwpos37_45 in37_45 sp37_45 78000.000000
Rwpos37_46 in37_46 sp37_46 78000.000000
Rwpos37_47 in37_47 sp37_47 78000.000000
Rwpos37_48 in37_48 sp37_48 78000.000000
Rwpos37_49 in37_49 sp37_49 78000.000000
Rwpos37_50 in37_50 sp37_50 78000.000000
Rwpos37_51 in37_51 sp37_51 202000.000000
Rwpos37_52 in37_52 sp37_52 78000.000000
Rwpos37_53 in37_53 sp37_53 202000.000000
Rwpos37_54 in37_54 sp37_54 202000.000000
Rwpos37_55 in37_55 sp37_55 202000.000000
Rwpos37_56 in37_56 sp37_56 202000.000000
Rwpos37_57 in37_57 sp37_57 78000.000000
Rwpos37_58 in37_58 sp37_58 202000.000000
Rwpos37_59 in37_59 sp37_59 78000.000000
Rwpos37_60 in37_60 sp37_60 202000.000000
Rwpos37_61 in37_61 sp37_61 78000.000000
Rwpos37_62 in37_62 sp37_62 202000.000000
Rwpos37_63 in37_63 sp37_63 202000.000000
Rwpos37_64 in37_64 sp37_64 202000.000000
Rwpos37_65 in37_65 sp37_65 78000.000000
Rwpos37_66 in37_66 sp37_66 202000.000000
Rwpos37_67 in37_67 sp37_67 78000.000000
Rwpos37_68 in37_68 sp37_68 202000.000000
Rwpos37_69 in37_69 sp37_69 202000.000000
Rwpos37_70 in37_70 sp37_70 78000.000000
Rwpos37_71 in37_71 sp37_71 202000.000000
Rwpos37_72 in37_72 sp37_72 78000.000000
Rwpos37_73 in37_73 sp37_73 78000.000000
Rwpos37_74 in37_74 sp37_74 78000.000000
Rwpos37_75 in37_75 sp37_75 78000.000000
Rwpos37_76 in37_76 sp37_76 78000.000000
Rwpos37_77 in37_77 sp37_77 78000.000000
Rwpos37_78 in37_78 sp37_78 78000.000000
Rwpos37_79 in37_79 sp37_79 202000.000000
Rwpos37_80 in37_80 sp37_80 202000.000000
Rwpos37_81 in37_81 sp37_81 202000.000000
Rwpos37_82 in37_82 sp37_82 202000.000000
Rwpos37_83 in37_83 sp37_83 202000.000000
Rwpos37_84 in37_84 sp37_84 202000.000000
Rwpos38_1 in38_1 sp38_1 78000.000000
Rwpos38_2 in38_2 sp38_2 202000.000000
Rwpos38_3 in38_3 sp38_3 202000.000000
Rwpos38_4 in38_4 sp38_4 202000.000000
Rwpos38_5 in38_5 sp38_5 202000.000000
Rwpos38_6 in38_6 sp38_6 78000.000000
Rwpos38_7 in38_7 sp38_7 202000.000000
Rwpos38_8 in38_8 sp38_8 202000.000000
Rwpos38_9 in38_9 sp38_9 202000.000000
Rwpos38_10 in38_10 sp38_10 202000.000000
Rwpos38_11 in38_11 sp38_11 78000.000000
Rwpos38_12 in38_12 sp38_12 202000.000000
Rwpos38_13 in38_13 sp38_13 78000.000000
Rwpos38_14 in38_14 sp38_14 202000.000000
Rwpos38_15 in38_15 sp38_15 78000.000000
Rwpos38_16 in38_16 sp38_16 202000.000000
Rwpos38_17 in38_17 sp38_17 78000.000000
Rwpos38_18 in38_18 sp38_18 202000.000000
Rwpos38_19 in38_19 sp38_19 202000.000000
Rwpos38_20 in38_20 sp38_20 78000.000000
Rwpos38_21 in38_21 sp38_21 78000.000000
Rwpos38_22 in38_22 sp38_22 78000.000000
Rwpos38_23 in38_23 sp38_23 78000.000000
Rwpos38_24 in38_24 sp38_24 78000.000000
Rwpos38_25 in38_25 sp38_25 78000.000000
Rwpos38_26 in38_26 sp38_26 78000.000000
Rwpos38_27 in38_27 sp38_27 202000.000000
Rwpos38_28 in38_28 sp38_28 202000.000000
Rwpos38_29 in38_29 sp38_29 202000.000000
Rwpos38_30 in38_30 sp38_30 202000.000000
Rwpos38_31 in38_31 sp38_31 78000.000000
Rwpos38_32 in38_32 sp38_32 78000.000000
Rwpos38_33 in38_33 sp38_33 78000.000000
Rwpos38_34 in38_34 sp38_34 202000.000000
Rwpos38_35 in38_35 sp38_35 202000.000000
Rwpos38_36 in38_36 sp38_36 202000.000000
Rwpos38_37 in38_37 sp38_37 78000.000000
Rwpos38_38 in38_38 sp38_38 202000.000000
Rwpos38_39 in38_39 sp38_39 202000.000000
Rwpos38_40 in38_40 sp38_40 78000.000000
Rwpos38_41 in38_41 sp38_41 202000.000000
Rwpos38_42 in38_42 sp38_42 78000.000000
Rwpos38_43 in38_43 sp38_43 78000.000000
Rwpos38_44 in38_44 sp38_44 78000.000000
Rwpos38_45 in38_45 sp38_45 202000.000000
Rwpos38_46 in38_46 sp38_46 202000.000000
Rwpos38_47 in38_47 sp38_47 202000.000000
Rwpos38_48 in38_48 sp38_48 202000.000000
Rwpos38_49 in38_49 sp38_49 202000.000000
Rwpos38_50 in38_50 sp38_50 202000.000000
Rwpos38_51 in38_51 sp38_51 78000.000000
Rwpos38_52 in38_52 sp38_52 202000.000000
Rwpos38_53 in38_53 sp38_53 202000.000000
Rwpos38_54 in38_54 sp38_54 78000.000000
Rwpos38_55 in38_55 sp38_55 202000.000000
Rwpos38_56 in38_56 sp38_56 78000.000000
Rwpos38_57 in38_57 sp38_57 78000.000000
Rwpos38_58 in38_58 sp38_58 78000.000000
Rwpos38_59 in38_59 sp38_59 202000.000000
Rwpos38_60 in38_60 sp38_60 202000.000000
Rwpos38_61 in38_61 sp38_61 202000.000000
Rwpos38_62 in38_62 sp38_62 78000.000000
Rwpos38_63 in38_63 sp38_63 202000.000000
Rwpos38_64 in38_64 sp38_64 78000.000000
Rwpos38_65 in38_65 sp38_65 202000.000000
Rwpos38_66 in38_66 sp38_66 202000.000000
Rwpos38_67 in38_67 sp38_67 202000.000000
Rwpos38_68 in38_68 sp38_68 78000.000000
Rwpos38_69 in38_69 sp38_69 202000.000000
Rwpos38_70 in38_70 sp38_70 78000.000000
Rwpos38_71 in38_71 sp38_71 202000.000000
Rwpos38_72 in38_72 sp38_72 78000.000000
Rwpos38_73 in38_73 sp38_73 78000.000000
Rwpos38_74 in38_74 sp38_74 202000.000000
Rwpos38_75 in38_75 sp38_75 202000.000000
Rwpos38_76 in38_76 sp38_76 202000.000000
Rwpos38_77 in38_77 sp38_77 202000.000000
Rwpos38_78 in38_78 sp38_78 202000.000000
Rwpos38_79 in38_79 sp38_79 202000.000000
Rwpos38_80 in38_80 sp38_80 78000.000000
Rwpos38_81 in38_81 sp38_81 78000.000000
Rwpos38_82 in38_82 sp38_82 202000.000000
Rwpos38_83 in38_83 sp38_83 202000.000000
Rwpos38_84 in38_84 sp38_84 202000.000000
Rwpos39_1 in39_1 sp39_1 78000.000000
Rwpos39_2 in39_2 sp39_2 78000.000000
Rwpos39_3 in39_3 sp39_3 78000.000000
Rwpos39_4 in39_4 sp39_4 78000.000000
Rwpos39_5 in39_5 sp39_5 78000.000000
Rwpos39_6 in39_6 sp39_6 78000.000000
Rwpos39_7 in39_7 sp39_7 202000.000000
Rwpos39_8 in39_8 sp39_8 78000.000000
Rwpos39_9 in39_9 sp39_9 78000.000000
Rwpos39_10 in39_10 sp39_10 202000.000000
Rwpos39_11 in39_11 sp39_11 202000.000000
Rwpos39_12 in39_12 sp39_12 202000.000000
Rwpos39_13 in39_13 sp39_13 78000.000000
Rwpos39_14 in39_14 sp39_14 78000.000000
Rwpos39_15 in39_15 sp39_15 202000.000000
Rwpos39_16 in39_16 sp39_16 78000.000000
Rwpos39_17 in39_17 sp39_17 202000.000000
Rwpos39_18 in39_18 sp39_18 78000.000000
Rwpos39_19 in39_19 sp39_19 202000.000000
Rwpos39_20 in39_20 sp39_20 78000.000000
Rwpos39_21 in39_21 sp39_21 202000.000000
Rwpos39_22 in39_22 sp39_22 202000.000000
Rwpos39_23 in39_23 sp39_23 78000.000000
Rwpos39_24 in39_24 sp39_24 202000.000000
Rwpos39_25 in39_25 sp39_25 78000.000000
Rwpos39_26 in39_26 sp39_26 78000.000000
Rwpos39_27 in39_27 sp39_27 78000.000000
Rwpos39_28 in39_28 sp39_28 202000.000000
Rwpos39_29 in39_29 sp39_29 78000.000000
Rwpos39_30 in39_30 sp39_30 78000.000000
Rwpos39_31 in39_31 sp39_31 202000.000000
Rwpos39_32 in39_32 sp39_32 78000.000000
Rwpos39_33 in39_33 sp39_33 202000.000000
Rwpos39_34 in39_34 sp39_34 202000.000000
Rwpos39_35 in39_35 sp39_35 78000.000000
Rwpos39_36 in39_36 sp39_36 202000.000000
Rwpos39_37 in39_37 sp39_37 202000.000000
Rwpos39_38 in39_38 sp39_38 202000.000000
Rwpos39_39 in39_39 sp39_39 78000.000000
Rwpos39_40 in39_40 sp39_40 202000.000000
Rwpos39_41 in39_41 sp39_41 78000.000000
Rwpos39_42 in39_42 sp39_42 78000.000000
Rwpos39_43 in39_43 sp39_43 202000.000000
Rwpos39_44 in39_44 sp39_44 78000.000000
Rwpos39_45 in39_45 sp39_45 78000.000000
Rwpos39_46 in39_46 sp39_46 78000.000000
Rwpos39_47 in39_47 sp39_47 78000.000000
Rwpos39_48 in39_48 sp39_48 202000.000000
Rwpos39_49 in39_49 sp39_49 202000.000000
Rwpos39_50 in39_50 sp39_50 202000.000000
Rwpos39_51 in39_51 sp39_51 202000.000000
Rwpos39_52 in39_52 sp39_52 202000.000000
Rwpos39_53 in39_53 sp39_53 78000.000000
Rwpos39_54 in39_54 sp39_54 78000.000000
Rwpos39_55 in39_55 sp39_55 202000.000000
Rwpos39_56 in39_56 sp39_56 78000.000000
Rwpos39_57 in39_57 sp39_57 202000.000000
Rwpos39_58 in39_58 sp39_58 78000.000000
Rwpos39_59 in39_59 sp39_59 78000.000000
Rwpos39_60 in39_60 sp39_60 78000.000000
Rwpos39_61 in39_61 sp39_61 202000.000000
Rwpos39_62 in39_62 sp39_62 202000.000000
Rwpos39_63 in39_63 sp39_63 202000.000000
Rwpos39_64 in39_64 sp39_64 202000.000000
Rwpos39_65 in39_65 sp39_65 202000.000000
Rwpos39_66 in39_66 sp39_66 78000.000000
Rwpos39_67 in39_67 sp39_67 202000.000000
Rwpos39_68 in39_68 sp39_68 202000.000000
Rwpos39_69 in39_69 sp39_69 202000.000000
Rwpos39_70 in39_70 sp39_70 202000.000000
Rwpos39_71 in39_71 sp39_71 78000.000000
Rwpos39_72 in39_72 sp39_72 78000.000000
Rwpos39_73 in39_73 sp39_73 202000.000000
Rwpos39_74 in39_74 sp39_74 78000.000000
Rwpos39_75 in39_75 sp39_75 78000.000000
Rwpos39_76 in39_76 sp39_76 78000.000000
Rwpos39_77 in39_77 sp39_77 78000.000000
Rwpos39_78 in39_78 sp39_78 78000.000000
Rwpos39_79 in39_79 sp39_79 78000.000000
Rwpos39_80 in39_80 sp39_80 78000.000000
Rwpos39_81 in39_81 sp39_81 78000.000000
Rwpos39_82 in39_82 sp39_82 202000.000000
Rwpos39_83 in39_83 sp39_83 78000.000000
Rwpos39_84 in39_84 sp39_84 78000.000000
Rwpos40_1 in40_1 sp40_1 78000.000000
Rwpos40_2 in40_2 sp40_2 202000.000000
Rwpos40_3 in40_3 sp40_3 202000.000000
Rwpos40_4 in40_4 sp40_4 202000.000000
Rwpos40_5 in40_5 sp40_5 202000.000000
Rwpos40_6 in40_6 sp40_6 202000.000000
Rwpos40_7 in40_7 sp40_7 78000.000000
Rwpos40_8 in40_8 sp40_8 202000.000000
Rwpos40_9 in40_9 sp40_9 202000.000000
Rwpos40_10 in40_10 sp40_10 202000.000000
Rwpos40_11 in40_11 sp40_11 78000.000000
Rwpos40_12 in40_12 sp40_12 202000.000000
Rwpos40_13 in40_13 sp40_13 78000.000000
Rwpos40_14 in40_14 sp40_14 202000.000000
Rwpos40_15 in40_15 sp40_15 202000.000000
Rwpos40_16 in40_16 sp40_16 78000.000000
Rwpos40_17 in40_17 sp40_17 78000.000000
Rwpos40_18 in40_18 sp40_18 202000.000000
Rwpos40_19 in40_19 sp40_19 78000.000000
Rwpos40_20 in40_20 sp40_20 78000.000000
Rwpos40_21 in40_21 sp40_21 78000.000000
Rwpos40_22 in40_22 sp40_22 78000.000000
Rwpos40_23 in40_23 sp40_23 202000.000000
Rwpos40_24 in40_24 sp40_24 78000.000000
Rwpos40_25 in40_25 sp40_25 78000.000000
Rwpos40_26 in40_26 sp40_26 78000.000000
Rwpos40_27 in40_27 sp40_27 202000.000000
Rwpos40_28 in40_28 sp40_28 78000.000000
Rwpos40_29 in40_29 sp40_29 78000.000000
Rwpos40_30 in40_30 sp40_30 78000.000000
Rwpos40_31 in40_31 sp40_31 202000.000000
Rwpos40_32 in40_32 sp40_32 78000.000000
Rwpos40_33 in40_33 sp40_33 78000.000000
Rwpos40_34 in40_34 sp40_34 202000.000000
Rwpos40_35 in40_35 sp40_35 202000.000000
Rwpos40_36 in40_36 sp40_36 78000.000000
Rwpos40_37 in40_37 sp40_37 78000.000000
Rwpos40_38 in40_38 sp40_38 202000.000000
Rwpos40_39 in40_39 sp40_39 78000.000000
Rwpos40_40 in40_40 sp40_40 78000.000000
Rwpos40_41 in40_41 sp40_41 78000.000000
Rwpos40_42 in40_42 sp40_42 202000.000000
Rwpos40_43 in40_43 sp40_43 78000.000000
Rwpos40_44 in40_44 sp40_44 78000.000000
Rwpos40_45 in40_45 sp40_45 202000.000000
Rwpos40_46 in40_46 sp40_46 202000.000000
Rwpos40_47 in40_47 sp40_47 78000.000000
Rwpos40_48 in40_48 sp40_48 78000.000000
Rwpos40_49 in40_49 sp40_49 202000.000000
Rwpos40_50 in40_50 sp40_50 78000.000000
Rwpos40_51 in40_51 sp40_51 78000.000000
Rwpos40_52 in40_52 sp40_52 202000.000000
Rwpos40_53 in40_53 sp40_53 202000.000000
Rwpos40_54 in40_54 sp40_54 202000.000000
Rwpos40_55 in40_55 sp40_55 78000.000000
Rwpos40_56 in40_56 sp40_56 202000.000000
Rwpos40_57 in40_57 sp40_57 78000.000000
Rwpos40_58 in40_58 sp40_58 202000.000000
Rwpos40_59 in40_59 sp40_59 78000.000000
Rwpos40_60 in40_60 sp40_60 78000.000000
Rwpos40_61 in40_61 sp40_61 78000.000000
Rwpos40_62 in40_62 sp40_62 78000.000000
Rwpos40_63 in40_63 sp40_63 78000.000000
Rwpos40_64 in40_64 sp40_64 202000.000000
Rwpos40_65 in40_65 sp40_65 202000.000000
Rwpos40_66 in40_66 sp40_66 78000.000000
Rwpos40_67 in40_67 sp40_67 78000.000000
Rwpos40_68 in40_68 sp40_68 78000.000000
Rwpos40_69 in40_69 sp40_69 202000.000000
Rwpos40_70 in40_70 sp40_70 78000.000000
Rwpos40_71 in40_71 sp40_71 78000.000000
Rwpos40_72 in40_72 sp40_72 202000.000000
Rwpos40_73 in40_73 sp40_73 202000.000000
Rwpos40_74 in40_74 sp40_74 202000.000000
Rwpos40_75 in40_75 sp40_75 78000.000000
Rwpos40_76 in40_76 sp40_76 78000.000000
Rwpos40_77 in40_77 sp40_77 202000.000000
Rwpos40_78 in40_78 sp40_78 78000.000000
Rwpos40_79 in40_79 sp40_79 78000.000000
Rwpos40_80 in40_80 sp40_80 202000.000000
Rwpos40_81 in40_81 sp40_81 78000.000000
Rwpos40_82 in40_82 sp40_82 202000.000000
Rwpos40_83 in40_83 sp40_83 202000.000000
Rwpos40_84 in40_84 sp40_84 202000.000000
Rwpos41_1 in41_1 sp41_1 78000.000000
Rwpos41_2 in41_2 sp41_2 202000.000000
Rwpos41_3 in41_3 sp41_3 202000.000000
Rwpos41_4 in41_4 sp41_4 78000.000000
Rwpos41_5 in41_5 sp41_5 202000.000000
Rwpos41_6 in41_6 sp41_6 78000.000000
Rwpos41_7 in41_7 sp41_7 202000.000000
Rwpos41_8 in41_8 sp41_8 78000.000000
Rwpos41_9 in41_9 sp41_9 78000.000000
Rwpos41_10 in41_10 sp41_10 78000.000000
Rwpos41_11 in41_11 sp41_11 78000.000000
Rwpos41_12 in41_12 sp41_12 202000.000000
Rwpos41_13 in41_13 sp41_13 78000.000000
Rwpos41_14 in41_14 sp41_14 202000.000000
Rwpos41_15 in41_15 sp41_15 202000.000000
Rwpos41_16 in41_16 sp41_16 202000.000000
Rwpos41_17 in41_17 sp41_17 78000.000000
Rwpos41_18 in41_18 sp41_18 78000.000000
Rwpos41_19 in41_19 sp41_19 202000.000000
Rwpos41_20 in41_20 sp41_20 78000.000000
Rwpos41_21 in41_21 sp41_21 78000.000000
Rwpos41_22 in41_22 sp41_22 78000.000000
Rwpos41_23 in41_23 sp41_23 78000.000000
Rwpos41_24 in41_24 sp41_24 78000.000000
Rwpos41_25 in41_25 sp41_25 78000.000000
Rwpos41_26 in41_26 sp41_26 78000.000000
Rwpos41_27 in41_27 sp41_27 202000.000000
Rwpos41_28 in41_28 sp41_28 202000.000000
Rwpos41_29 in41_29 sp41_29 202000.000000
Rwpos41_30 in41_30 sp41_30 202000.000000
Rwpos41_31 in41_31 sp41_31 202000.000000
Rwpos41_32 in41_32 sp41_32 202000.000000
Rwpos41_33 in41_33 sp41_33 202000.000000
Rwpos41_34 in41_34 sp41_34 78000.000000
Rwpos41_35 in41_35 sp41_35 202000.000000
Rwpos41_36 in41_36 sp41_36 78000.000000
Rwpos41_37 in41_37 sp41_37 202000.000000
Rwpos41_38 in41_38 sp41_38 202000.000000
Rwpos41_39 in41_39 sp41_39 78000.000000
Rwpos41_40 in41_40 sp41_40 78000.000000
Rwpos41_41 in41_41 sp41_41 78000.000000
Rwpos41_42 in41_42 sp41_42 78000.000000
Rwpos41_43 in41_43 sp41_43 78000.000000
Rwpos41_44 in41_44 sp41_44 78000.000000
Rwpos41_45 in41_45 sp41_45 78000.000000
Rwpos41_46 in41_46 sp41_46 78000.000000
Rwpos41_47 in41_47 sp41_47 78000.000000
Rwpos41_48 in41_48 sp41_48 202000.000000
Rwpos41_49 in41_49 sp41_49 202000.000000
Rwpos41_50 in41_50 sp41_50 202000.000000
Rwpos41_51 in41_51 sp41_51 202000.000000
Rwpos41_52 in41_52 sp41_52 202000.000000
Rwpos41_53 in41_53 sp41_53 202000.000000
Rwpos41_54 in41_54 sp41_54 202000.000000
Rwpos41_55 in41_55 sp41_55 202000.000000
Rwpos41_56 in41_56 sp41_56 78000.000000
Rwpos41_57 in41_57 sp41_57 78000.000000
Rwpos41_58 in41_58 sp41_58 78000.000000
Rwpos41_59 in41_59 sp41_59 78000.000000
Rwpos41_60 in41_60 sp41_60 78000.000000
Rwpos41_61 in41_61 sp41_61 202000.000000
Rwpos41_62 in41_62 sp41_62 78000.000000
Rwpos41_63 in41_63 sp41_63 202000.000000
Rwpos41_64 in41_64 sp41_64 78000.000000
Rwpos41_65 in41_65 sp41_65 78000.000000
Rwpos41_66 in41_66 sp41_66 202000.000000
Rwpos41_67 in41_67 sp41_67 78000.000000
Rwpos41_68 in41_68 sp41_68 78000.000000
Rwpos41_69 in41_69 sp41_69 202000.000000
Rwpos41_70 in41_70 sp41_70 78000.000000
Rwpos41_71 in41_71 sp41_71 78000.000000
Rwpos41_72 in41_72 sp41_72 202000.000000
Rwpos41_73 in41_73 sp41_73 202000.000000
Rwpos41_74 in41_74 sp41_74 202000.000000
Rwpos41_75 in41_75 sp41_75 78000.000000
Rwpos41_76 in41_76 sp41_76 202000.000000
Rwpos41_77 in41_77 sp41_77 78000.000000
Rwpos41_78 in41_78 sp41_78 202000.000000
Rwpos41_79 in41_79 sp41_79 202000.000000
Rwpos41_80 in41_80 sp41_80 78000.000000
Rwpos41_81 in41_81 sp41_81 78000.000000
Rwpos41_82 in41_82 sp41_82 202000.000000
Rwpos41_83 in41_83 sp41_83 78000.000000
Rwpos41_84 in41_84 sp41_84 78000.000000
Rwpos42_1 in42_1 sp42_1 78000.000000
Rwpos42_2 in42_2 sp42_2 202000.000000
Rwpos42_3 in42_3 sp42_3 78000.000000
Rwpos42_4 in42_4 sp42_4 78000.000000
Rwpos42_5 in42_5 sp42_5 78000.000000
Rwpos42_6 in42_6 sp42_6 78000.000000
Rwpos42_7 in42_7 sp42_7 78000.000000
Rwpos42_8 in42_8 sp42_8 78000.000000
Rwpos42_9 in42_9 sp42_9 78000.000000
Rwpos42_10 in42_10 sp42_10 78000.000000
Rwpos42_11 in42_11 sp42_11 202000.000000
Rwpos42_12 in42_12 sp42_12 78000.000000
Rwpos42_13 in42_13 sp42_13 78000.000000
Rwpos42_14 in42_14 sp42_14 202000.000000
Rwpos42_15 in42_15 sp42_15 78000.000000
Rwpos42_16 in42_16 sp42_16 78000.000000
Rwpos42_17 in42_17 sp42_17 202000.000000
Rwpos42_18 in42_18 sp42_18 78000.000000
Rwpos42_19 in42_19 sp42_19 78000.000000
Rwpos42_20 in42_20 sp42_20 78000.000000
Rwpos42_21 in42_21 sp42_21 202000.000000
Rwpos42_22 in42_22 sp42_22 78000.000000
Rwpos42_23 in42_23 sp42_23 202000.000000
Rwpos42_24 in42_24 sp42_24 202000.000000
Rwpos42_25 in42_25 sp42_25 78000.000000
Rwpos42_26 in42_26 sp42_26 78000.000000
Rwpos42_27 in42_27 sp42_27 78000.000000
Rwpos42_28 in42_28 sp42_28 78000.000000
Rwpos42_29 in42_29 sp42_29 202000.000000
Rwpos42_30 in42_30 sp42_30 78000.000000
Rwpos42_31 in42_31 sp42_31 202000.000000
Rwpos42_32 in42_32 sp42_32 202000.000000
Rwpos42_33 in42_33 sp42_33 78000.000000
Rwpos42_34 in42_34 sp42_34 78000.000000
Rwpos42_35 in42_35 sp42_35 78000.000000
Rwpos42_36 in42_36 sp42_36 78000.000000
Rwpos42_37 in42_37 sp42_37 202000.000000
Rwpos42_38 in42_38 sp42_38 78000.000000
Rwpos42_39 in42_39 sp42_39 78000.000000
Rwpos42_40 in42_40 sp42_40 202000.000000
Rwpos42_41 in42_41 sp42_41 202000.000000
Rwpos42_42 in42_42 sp42_42 202000.000000
Rwpos42_43 in42_43 sp42_43 78000.000000
Rwpos42_44 in42_44 sp42_44 202000.000000
Rwpos42_45 in42_45 sp42_45 78000.000000
Rwpos42_46 in42_46 sp42_46 202000.000000
Rwpos42_47 in42_47 sp42_47 78000.000000
Rwpos42_48 in42_48 sp42_48 202000.000000
Rwpos42_49 in42_49 sp42_49 202000.000000
Rwpos42_50 in42_50 sp42_50 202000.000000
Rwpos42_51 in42_51 sp42_51 202000.000000
Rwpos42_52 in42_52 sp42_52 202000.000000
Rwpos42_53 in42_53 sp42_53 78000.000000
Rwpos42_54 in42_54 sp42_54 78000.000000
Rwpos42_55 in42_55 sp42_55 202000.000000
Rwpos42_56 in42_56 sp42_56 78000.000000
Rwpos42_57 in42_57 sp42_57 78000.000000
Rwpos42_58 in42_58 sp42_58 202000.000000
Rwpos42_59 in42_59 sp42_59 202000.000000
Rwpos42_60 in42_60 sp42_60 78000.000000
Rwpos42_61 in42_61 sp42_61 202000.000000
Rwpos42_62 in42_62 sp42_62 202000.000000
Rwpos42_63 in42_63 sp42_63 78000.000000
Rwpos42_64 in42_64 sp42_64 202000.000000
Rwpos42_65 in42_65 sp42_65 78000.000000
Rwpos42_66 in42_66 sp42_66 202000.000000
Rwpos42_67 in42_67 sp42_67 202000.000000
Rwpos42_68 in42_68 sp42_68 202000.000000
Rwpos42_69 in42_69 sp42_69 202000.000000
Rwpos42_70 in42_70 sp42_70 202000.000000
Rwpos42_71 in42_71 sp42_71 78000.000000
Rwpos42_72 in42_72 sp42_72 78000.000000
Rwpos42_73 in42_73 sp42_73 202000.000000
Rwpos42_74 in42_74 sp42_74 202000.000000
Rwpos42_75 in42_75 sp42_75 78000.000000
Rwpos42_76 in42_76 sp42_76 202000.000000
Rwpos42_77 in42_77 sp42_77 78000.000000
Rwpos42_78 in42_78 sp42_78 202000.000000
Rwpos42_79 in42_79 sp42_79 202000.000000
Rwpos42_80 in42_80 sp42_80 78000.000000
Rwpos42_81 in42_81 sp42_81 202000.000000
Rwpos42_82 in42_82 sp42_82 78000.000000
Rwpos42_83 in42_83 sp42_83 78000.000000
Rwpos42_84 in42_84 sp42_84 78000.000000
Rwpos43_1 in43_1 sp43_1 78000.000000
Rwpos43_2 in43_2 sp43_2 202000.000000
Rwpos43_3 in43_3 sp43_3 202000.000000
Rwpos43_4 in43_4 sp43_4 78000.000000
Rwpos43_5 in43_5 sp43_5 78000.000000
Rwpos43_6 in43_6 sp43_6 202000.000000
Rwpos43_7 in43_7 sp43_7 78000.000000
Rwpos43_8 in43_8 sp43_8 78000.000000
Rwpos43_9 in43_9 sp43_9 78000.000000
Rwpos43_10 in43_10 sp43_10 78000.000000
Rwpos43_11 in43_11 sp43_11 202000.000000
Rwpos43_12 in43_12 sp43_12 202000.000000
Rwpos43_13 in43_13 sp43_13 78000.000000
Rwpos43_14 in43_14 sp43_14 78000.000000
Rwpos43_15 in43_15 sp43_15 202000.000000
Rwpos43_16 in43_16 sp43_16 78000.000000
Rwpos43_17 in43_17 sp43_17 202000.000000
Rwpos43_18 in43_18 sp43_18 202000.000000
Rwpos43_19 in43_19 sp43_19 78000.000000
Rwpos43_20 in43_20 sp43_20 78000.000000
Rwpos43_21 in43_21 sp43_21 202000.000000
Rwpos43_22 in43_22 sp43_22 78000.000000
Rwpos43_23 in43_23 sp43_23 202000.000000
Rwpos43_24 in43_24 sp43_24 202000.000000
Rwpos43_25 in43_25 sp43_25 202000.000000
Rwpos43_26 in43_26 sp43_26 78000.000000
Rwpos43_27 in43_27 sp43_27 78000.000000
Rwpos43_28 in43_28 sp43_28 78000.000000
Rwpos43_29 in43_29 sp43_29 78000.000000
Rwpos43_30 in43_30 sp43_30 202000.000000
Rwpos43_31 in43_31 sp43_31 78000.000000
Rwpos43_32 in43_32 sp43_32 78000.000000
Rwpos43_33 in43_33 sp43_33 202000.000000
Rwpos43_34 in43_34 sp43_34 78000.000000
Rwpos43_35 in43_35 sp43_35 202000.000000
Rwpos43_36 in43_36 sp43_36 78000.000000
Rwpos43_37 in43_37 sp43_37 78000.000000
Rwpos43_38 in43_38 sp43_38 78000.000000
Rwpos43_39 in43_39 sp43_39 78000.000000
Rwpos43_40 in43_40 sp43_40 78000.000000
Rwpos43_41 in43_41 sp43_41 78000.000000
Rwpos43_42 in43_42 sp43_42 202000.000000
Rwpos43_43 in43_43 sp43_43 202000.000000
Rwpos43_44 in43_44 sp43_44 202000.000000
Rwpos43_45 in43_45 sp43_45 78000.000000
Rwpos43_46 in43_46 sp43_46 78000.000000
Rwpos43_47 in43_47 sp43_47 202000.000000
Rwpos43_48 in43_48 sp43_48 202000.000000
Rwpos43_49 in43_49 sp43_49 78000.000000
Rwpos43_50 in43_50 sp43_50 78000.000000
Rwpos43_51 in43_51 sp43_51 202000.000000
Rwpos43_52 in43_52 sp43_52 78000.000000
Rwpos43_53 in43_53 sp43_53 78000.000000
Rwpos43_54 in43_54 sp43_54 78000.000000
Rwpos43_55 in43_55 sp43_55 78000.000000
Rwpos43_56 in43_56 sp43_56 78000.000000
Rwpos43_57 in43_57 sp43_57 202000.000000
Rwpos43_58 in43_58 sp43_58 78000.000000
Rwpos43_59 in43_59 sp43_59 202000.000000
Rwpos43_60 in43_60 sp43_60 78000.000000
Rwpos43_61 in43_61 sp43_61 78000.000000
Rwpos43_62 in43_62 sp43_62 202000.000000
Rwpos43_63 in43_63 sp43_63 78000.000000
Rwpos43_64 in43_64 sp43_64 202000.000000
Rwpos43_65 in43_65 sp43_65 202000.000000
Rwpos43_66 in43_66 sp43_66 78000.000000
Rwpos43_67 in43_67 sp43_67 78000.000000
Rwpos43_68 in43_68 sp43_68 202000.000000
Rwpos43_69 in43_69 sp43_69 78000.000000
Rwpos43_70 in43_70 sp43_70 78000.000000
Rwpos43_71 in43_71 sp43_71 78000.000000
Rwpos43_72 in43_72 sp43_72 202000.000000
Rwpos43_73 in43_73 sp43_73 78000.000000
Rwpos43_74 in43_74 sp43_74 78000.000000
Rwpos43_75 in43_75 sp43_75 78000.000000
Rwpos43_76 in43_76 sp43_76 78000.000000
Rwpos43_77 in43_77 sp43_77 202000.000000
Rwpos43_78 in43_78 sp43_78 202000.000000
Rwpos43_79 in43_79 sp43_79 78000.000000
Rwpos43_80 in43_80 sp43_80 202000.000000
Rwpos43_81 in43_81 sp43_81 202000.000000
Rwpos43_82 in43_82 sp43_82 78000.000000
Rwpos43_83 in43_83 sp43_83 202000.000000
Rwpos43_84 in43_84 sp43_84 202000.000000
Rwpos44_1 in44_1 sp44_1 202000.000000
Rwpos44_2 in44_2 sp44_2 202000.000000
Rwpos44_3 in44_3 sp44_3 78000.000000
Rwpos44_4 in44_4 sp44_4 202000.000000
Rwpos44_5 in44_5 sp44_5 78000.000000
Rwpos44_6 in44_6 sp44_6 202000.000000
Rwpos44_7 in44_7 sp44_7 202000.000000
Rwpos44_8 in44_8 sp44_8 78000.000000
Rwpos44_9 in44_9 sp44_9 78000.000000
Rwpos44_10 in44_10 sp44_10 78000.000000
Rwpos44_11 in44_11 sp44_11 202000.000000
Rwpos44_12 in44_12 sp44_12 202000.000000
Rwpos44_13 in44_13 sp44_13 78000.000000
Rwpos44_14 in44_14 sp44_14 78000.000000
Rwpos44_15 in44_15 sp44_15 202000.000000
Rwpos44_16 in44_16 sp44_16 202000.000000
Rwpos44_17 in44_17 sp44_17 202000.000000
Rwpos44_18 in44_18 sp44_18 78000.000000
Rwpos44_19 in44_19 sp44_19 78000.000000
Rwpos44_20 in44_20 sp44_20 78000.000000
Rwpos44_21 in44_21 sp44_21 78000.000000
Rwpos44_22 in44_22 sp44_22 78000.000000
Rwpos44_23 in44_23 sp44_23 202000.000000
Rwpos44_24 in44_24 sp44_24 202000.000000
Rwpos44_25 in44_25 sp44_25 78000.000000
Rwpos44_26 in44_26 sp44_26 78000.000000
Rwpos44_27 in44_27 sp44_27 78000.000000
Rwpos44_28 in44_28 sp44_28 202000.000000
Rwpos44_29 in44_29 sp44_29 78000.000000
Rwpos44_30 in44_30 sp44_30 78000.000000
Rwpos44_31 in44_31 sp44_31 78000.000000
Rwpos44_32 in44_32 sp44_32 202000.000000
Rwpos44_33 in44_33 sp44_33 78000.000000
Rwpos44_34 in44_34 sp44_34 78000.000000
Rwpos44_35 in44_35 sp44_35 78000.000000
Rwpos44_36 in44_36 sp44_36 202000.000000
Rwpos44_37 in44_37 sp44_37 202000.000000
Rwpos44_38 in44_38 sp44_38 78000.000000
Rwpos44_39 in44_39 sp44_39 78000.000000
Rwpos44_40 in44_40 sp44_40 202000.000000
Rwpos44_41 in44_41 sp44_41 202000.000000
Rwpos44_42 in44_42 sp44_42 202000.000000
Rwpos44_43 in44_43 sp44_43 78000.000000
Rwpos44_44 in44_44 sp44_44 202000.000000
Rwpos44_45 in44_45 sp44_45 78000.000000
Rwpos44_46 in44_46 sp44_46 78000.000000
Rwpos44_47 in44_47 sp44_47 78000.000000
Rwpos44_48 in44_48 sp44_48 202000.000000
Rwpos44_49 in44_49 sp44_49 78000.000000
Rwpos44_50 in44_50 sp44_50 78000.000000
Rwpos44_51 in44_51 sp44_51 78000.000000
Rwpos44_52 in44_52 sp44_52 78000.000000
Rwpos44_53 in44_53 sp44_53 202000.000000
Rwpos44_54 in44_54 sp44_54 78000.000000
Rwpos44_55 in44_55 sp44_55 78000.000000
Rwpos44_56 in44_56 sp44_56 202000.000000
Rwpos44_57 in44_57 sp44_57 202000.000000
Rwpos44_58 in44_58 sp44_58 78000.000000
Rwpos44_59 in44_59 sp44_59 202000.000000
Rwpos44_60 in44_60 sp44_60 202000.000000
Rwpos44_61 in44_61 sp44_61 202000.000000
Rwpos44_62 in44_62 sp44_62 202000.000000
Rwpos44_63 in44_63 sp44_63 78000.000000
Rwpos44_64 in44_64 sp44_64 202000.000000
Rwpos44_65 in44_65 sp44_65 202000.000000
Rwpos44_66 in44_66 sp44_66 78000.000000
Rwpos44_67 in44_67 sp44_67 78000.000000
Rwpos44_68 in44_68 sp44_68 202000.000000
Rwpos44_69 in44_69 sp44_69 78000.000000
Rwpos44_70 in44_70 sp44_70 78000.000000
Rwpos44_71 in44_71 sp44_71 78000.000000
Rwpos44_72 in44_72 sp44_72 78000.000000
Rwpos44_73 in44_73 sp44_73 202000.000000
Rwpos44_74 in44_74 sp44_74 202000.000000
Rwpos44_75 in44_75 sp44_75 78000.000000
Rwpos44_76 in44_76 sp44_76 78000.000000
Rwpos44_77 in44_77 sp44_77 78000.000000
Rwpos44_78 in44_78 sp44_78 202000.000000
Rwpos44_79 in44_79 sp44_79 202000.000000
Rwpos44_80 in44_80 sp44_80 78000.000000
Rwpos44_81 in44_81 sp44_81 202000.000000
Rwpos44_82 in44_82 sp44_82 78000.000000
Rwpos44_83 in44_83 sp44_83 202000.000000
Rwpos44_84 in44_84 sp44_84 78000.000000
Rwpos45_1 in45_1 sp45_1 202000.000000
Rwpos45_2 in45_2 sp45_2 202000.000000
Rwpos45_3 in45_3 sp45_3 78000.000000
Rwpos45_4 in45_4 sp45_4 202000.000000
Rwpos45_5 in45_5 sp45_5 78000.000000
Rwpos45_6 in45_6 sp45_6 202000.000000
Rwpos45_7 in45_7 sp45_7 202000.000000
Rwpos45_8 in45_8 sp45_8 202000.000000
Rwpos45_9 in45_9 sp45_9 202000.000000
Rwpos45_10 in45_10 sp45_10 78000.000000
Rwpos45_11 in45_11 sp45_11 78000.000000
Rwpos45_12 in45_12 sp45_12 202000.000000
Rwpos45_13 in45_13 sp45_13 202000.000000
Rwpos45_14 in45_14 sp45_14 202000.000000
Rwpos45_15 in45_15 sp45_15 78000.000000
Rwpos45_16 in45_16 sp45_16 202000.000000
Rwpos45_17 in45_17 sp45_17 202000.000000
Rwpos45_18 in45_18 sp45_18 78000.000000
Rwpos45_19 in45_19 sp45_19 78000.000000
Rwpos45_20 in45_20 sp45_20 78000.000000
Rwpos45_21 in45_21 sp45_21 202000.000000
Rwpos45_22 in45_22 sp45_22 202000.000000
Rwpos45_23 in45_23 sp45_23 78000.000000
Rwpos45_24 in45_24 sp45_24 202000.000000
Rwpos45_25 in45_25 sp45_25 78000.000000
Rwpos45_26 in45_26 sp45_26 202000.000000
Rwpos45_27 in45_27 sp45_27 202000.000000
Rwpos45_28 in45_28 sp45_28 202000.000000
Rwpos45_29 in45_29 sp45_29 202000.000000
Rwpos45_30 in45_30 sp45_30 202000.000000
Rwpos45_31 in45_31 sp45_31 202000.000000
Rwpos45_32 in45_32 sp45_32 78000.000000
Rwpos45_33 in45_33 sp45_33 78000.000000
Rwpos45_34 in45_34 sp45_34 202000.000000
Rwpos45_35 in45_35 sp45_35 78000.000000
Rwpos45_36 in45_36 sp45_36 202000.000000
Rwpos45_37 in45_37 sp45_37 202000.000000
Rwpos45_38 in45_38 sp45_38 202000.000000
Rwpos45_39 in45_39 sp45_39 202000.000000
Rwpos45_40 in45_40 sp45_40 78000.000000
Rwpos45_41 in45_41 sp45_41 78000.000000
Rwpos45_42 in45_42 sp45_42 202000.000000
Rwpos45_43 in45_43 sp45_43 202000.000000
Rwpos45_44 in45_44 sp45_44 78000.000000
Rwpos45_45 in45_45 sp45_45 78000.000000
Rwpos45_46 in45_46 sp45_46 202000.000000
Rwpos45_47 in45_47 sp45_47 202000.000000
Rwpos45_48 in45_48 sp45_48 78000.000000
Rwpos45_49 in45_49 sp45_49 78000.000000
Rwpos45_50 in45_50 sp45_50 78000.000000
Rwpos45_51 in45_51 sp45_51 202000.000000
Rwpos45_52 in45_52 sp45_52 202000.000000
Rwpos45_53 in45_53 sp45_53 202000.000000
Rwpos45_54 in45_54 sp45_54 202000.000000
Rwpos45_55 in45_55 sp45_55 78000.000000
Rwpos45_56 in45_56 sp45_56 78000.000000
Rwpos45_57 in45_57 sp45_57 78000.000000
Rwpos45_58 in45_58 sp45_58 78000.000000
Rwpos45_59 in45_59 sp45_59 202000.000000
Rwpos45_60 in45_60 sp45_60 202000.000000
Rwpos45_61 in45_61 sp45_61 78000.000000
Rwpos45_62 in45_62 sp45_62 202000.000000
Rwpos45_63 in45_63 sp45_63 78000.000000
Rwpos45_64 in45_64 sp45_64 202000.000000
Rwpos45_65 in45_65 sp45_65 78000.000000
Rwpos45_66 in45_66 sp45_66 78000.000000
Rwpos45_67 in45_67 sp45_67 202000.000000
Rwpos45_68 in45_68 sp45_68 202000.000000
Rwpos45_69 in45_69 sp45_69 78000.000000
Rwpos45_70 in45_70 sp45_70 202000.000000
Rwpos45_71 in45_71 sp45_71 78000.000000
Rwpos45_72 in45_72 sp45_72 202000.000000
Rwpos45_73 in45_73 sp45_73 202000.000000
Rwpos45_74 in45_74 sp45_74 78000.000000
Rwpos45_75 in45_75 sp45_75 78000.000000
Rwpos45_76 in45_76 sp45_76 202000.000000
Rwpos45_77 in45_77 sp45_77 78000.000000
Rwpos45_78 in45_78 sp45_78 202000.000000
Rwpos45_79 in45_79 sp45_79 78000.000000
Rwpos45_80 in45_80 sp45_80 78000.000000
Rwpos45_81 in45_81 sp45_81 78000.000000
Rwpos45_82 in45_82 sp45_82 202000.000000
Rwpos45_83 in45_83 sp45_83 78000.000000
Rwpos45_84 in45_84 sp45_84 78000.000000
Rwpos46_1 in46_1 sp46_1 78000.000000
Rwpos46_2 in46_2 sp46_2 78000.000000
Rwpos46_3 in46_3 sp46_3 78000.000000
Rwpos46_4 in46_4 sp46_4 202000.000000
Rwpos46_5 in46_5 sp46_5 78000.000000
Rwpos46_6 in46_6 sp46_6 78000.000000
Rwpos46_7 in46_7 sp46_7 78000.000000
Rwpos46_8 in46_8 sp46_8 202000.000000
Rwpos46_9 in46_9 sp46_9 202000.000000
Rwpos46_10 in46_10 sp46_10 202000.000000
Rwpos46_11 in46_11 sp46_11 78000.000000
Rwpos46_12 in46_12 sp46_12 202000.000000
Rwpos46_13 in46_13 sp46_13 78000.000000
Rwpos46_14 in46_14 sp46_14 78000.000000
Rwpos46_15 in46_15 sp46_15 78000.000000
Rwpos46_16 in46_16 sp46_16 202000.000000
Rwpos46_17 in46_17 sp46_17 78000.000000
Rwpos46_18 in46_18 sp46_18 78000.000000
Rwpos46_19 in46_19 sp46_19 202000.000000
Rwpos46_20 in46_20 sp46_20 202000.000000
Rwpos46_21 in46_21 sp46_21 202000.000000
Rwpos46_22 in46_22 sp46_22 78000.000000
Rwpos46_23 in46_23 sp46_23 78000.000000
Rwpos46_24 in46_24 sp46_24 78000.000000
Rwpos46_25 in46_25 sp46_25 78000.000000
Rwpos46_26 in46_26 sp46_26 78000.000000
Rwpos46_27 in46_27 sp46_27 202000.000000
Rwpos46_28 in46_28 sp46_28 202000.000000
Rwpos46_29 in46_29 sp46_29 202000.000000
Rwpos46_30 in46_30 sp46_30 202000.000000
Rwpos46_31 in46_31 sp46_31 78000.000000
Rwpos46_32 in46_32 sp46_32 78000.000000
Rwpos46_33 in46_33 sp46_33 78000.000000
Rwpos46_34 in46_34 sp46_34 202000.000000
Rwpos46_35 in46_35 sp46_35 78000.000000
Rwpos46_36 in46_36 sp46_36 78000.000000
Rwpos46_37 in46_37 sp46_37 202000.000000
Rwpos46_38 in46_38 sp46_38 78000.000000
Rwpos46_39 in46_39 sp46_39 78000.000000
Rwpos46_40 in46_40 sp46_40 202000.000000
Rwpos46_41 in46_41 sp46_41 78000.000000
Rwpos46_42 in46_42 sp46_42 78000.000000
Rwpos46_43 in46_43 sp46_43 202000.000000
Rwpos46_44 in46_44 sp46_44 202000.000000
Rwpos46_45 in46_45 sp46_45 202000.000000
Rwpos46_46 in46_46 sp46_46 78000.000000
Rwpos46_47 in46_47 sp46_47 78000.000000
Rwpos46_48 in46_48 sp46_48 202000.000000
Rwpos46_49 in46_49 sp46_49 202000.000000
Rwpos46_50 in46_50 sp46_50 202000.000000
Rwpos46_51 in46_51 sp46_51 78000.000000
Rwpos46_52 in46_52 sp46_52 202000.000000
Rwpos46_53 in46_53 sp46_53 202000.000000
Rwpos46_54 in46_54 sp46_54 202000.000000
Rwpos46_55 in46_55 sp46_55 202000.000000
Rwpos46_56 in46_56 sp46_56 78000.000000
Rwpos46_57 in46_57 sp46_57 78000.000000
Rwpos46_58 in46_58 sp46_58 78000.000000
Rwpos46_59 in46_59 sp46_59 78000.000000
Rwpos46_60 in46_60 sp46_60 202000.000000
Rwpos46_61 in46_61 sp46_61 78000.000000
Rwpos46_62 in46_62 sp46_62 78000.000000
Rwpos46_63 in46_63 sp46_63 202000.000000
Rwpos46_64 in46_64 sp46_64 202000.000000
Rwpos46_65 in46_65 sp46_65 78000.000000
Rwpos46_66 in46_66 sp46_66 202000.000000
Rwpos46_67 in46_67 sp46_67 78000.000000
Rwpos46_68 in46_68 sp46_68 202000.000000
Rwpos46_69 in46_69 sp46_69 202000.000000
Rwpos46_70 in46_70 sp46_70 78000.000000
Rwpos46_71 in46_71 sp46_71 202000.000000
Rwpos46_72 in46_72 sp46_72 78000.000000
Rwpos46_73 in46_73 sp46_73 202000.000000
Rwpos46_74 in46_74 sp46_74 78000.000000
Rwpos46_75 in46_75 sp46_75 78000.000000
Rwpos46_76 in46_76 sp46_76 78000.000000
Rwpos46_77 in46_77 sp46_77 78000.000000
Rwpos46_78 in46_78 sp46_78 202000.000000
Rwpos46_79 in46_79 sp46_79 78000.000000
Rwpos46_80 in46_80 sp46_80 78000.000000
Rwpos46_81 in46_81 sp46_81 78000.000000
Rwpos46_82 in46_82 sp46_82 202000.000000
Rwpos46_83 in46_83 sp46_83 78000.000000
Rwpos46_84 in46_84 sp46_84 78000.000000
Rwpos47_1 in47_1 sp47_1 78000.000000
Rwpos47_2 in47_2 sp47_2 78000.000000
Rwpos47_3 in47_3 sp47_3 202000.000000
Rwpos47_4 in47_4 sp47_4 202000.000000
Rwpos47_5 in47_5 sp47_5 202000.000000
Rwpos47_6 in47_6 sp47_6 202000.000000
Rwpos47_7 in47_7 sp47_7 78000.000000
Rwpos47_8 in47_8 sp47_8 78000.000000
Rwpos47_9 in47_9 sp47_9 78000.000000
Rwpos47_10 in47_10 sp47_10 78000.000000
Rwpos47_11 in47_11 sp47_11 78000.000000
Rwpos47_12 in47_12 sp47_12 78000.000000
Rwpos47_13 in47_13 sp47_13 202000.000000
Rwpos47_14 in47_14 sp47_14 78000.000000
Rwpos47_15 in47_15 sp47_15 78000.000000
Rwpos47_16 in47_16 sp47_16 78000.000000
Rwpos47_17 in47_17 sp47_17 202000.000000
Rwpos47_18 in47_18 sp47_18 78000.000000
Rwpos47_19 in47_19 sp47_19 78000.000000
Rwpos47_20 in47_20 sp47_20 78000.000000
Rwpos47_21 in47_21 sp47_21 78000.000000
Rwpos47_22 in47_22 sp47_22 202000.000000
Rwpos47_23 in47_23 sp47_23 78000.000000
Rwpos47_24 in47_24 sp47_24 202000.000000
Rwpos47_25 in47_25 sp47_25 202000.000000
Rwpos47_26 in47_26 sp47_26 78000.000000
Rwpos47_27 in47_27 sp47_27 202000.000000
Rwpos47_28 in47_28 sp47_28 78000.000000
Rwpos47_29 in47_29 sp47_29 202000.000000
Rwpos47_30 in47_30 sp47_30 202000.000000
Rwpos47_31 in47_31 sp47_31 202000.000000
Rwpos47_32 in47_32 sp47_32 78000.000000
Rwpos47_33 in47_33 sp47_33 78000.000000
Rwpos47_34 in47_34 sp47_34 78000.000000
Rwpos47_35 in47_35 sp47_35 202000.000000
Rwpos47_36 in47_36 sp47_36 78000.000000
Rwpos47_37 in47_37 sp47_37 78000.000000
Rwpos47_38 in47_38 sp47_38 78000.000000
Rwpos47_39 in47_39 sp47_39 202000.000000
Rwpos47_40 in47_40 sp47_40 78000.000000
Rwpos47_41 in47_41 sp47_41 202000.000000
Rwpos47_42 in47_42 sp47_42 78000.000000
Rwpos47_43 in47_43 sp47_43 78000.000000
Rwpos47_44 in47_44 sp47_44 78000.000000
Rwpos47_45 in47_45 sp47_45 78000.000000
Rwpos47_46 in47_46 sp47_46 202000.000000
Rwpos47_47 in47_47 sp47_47 202000.000000
Rwpos47_48 in47_48 sp47_48 78000.000000
Rwpos47_49 in47_49 sp47_49 78000.000000
Rwpos47_50 in47_50 sp47_50 78000.000000
Rwpos47_51 in47_51 sp47_51 78000.000000
Rwpos47_52 in47_52 sp47_52 78000.000000
Rwpos47_53 in47_53 sp47_53 202000.000000
Rwpos47_54 in47_54 sp47_54 202000.000000
Rwpos47_55 in47_55 sp47_55 202000.000000
Rwpos47_56 in47_56 sp47_56 78000.000000
Rwpos47_57 in47_57 sp47_57 202000.000000
Rwpos47_58 in47_58 sp47_58 78000.000000
Rwpos47_59 in47_59 sp47_59 78000.000000
Rwpos47_60 in47_60 sp47_60 78000.000000
Rwpos47_61 in47_61 sp47_61 78000.000000
Rwpos47_62 in47_62 sp47_62 202000.000000
Rwpos47_63 in47_63 sp47_63 78000.000000
Rwpos47_64 in47_64 sp47_64 202000.000000
Rwpos47_65 in47_65 sp47_65 202000.000000
Rwpos47_66 in47_66 sp47_66 78000.000000
Rwpos47_67 in47_67 sp47_67 78000.000000
Rwpos47_68 in47_68 sp47_68 202000.000000
Rwpos47_69 in47_69 sp47_69 78000.000000
Rwpos47_70 in47_70 sp47_70 202000.000000
Rwpos47_71 in47_71 sp47_71 78000.000000
Rwpos47_72 in47_72 sp47_72 78000.000000
Rwpos47_73 in47_73 sp47_73 78000.000000
Rwpos47_74 in47_74 sp47_74 202000.000000
Rwpos47_75 in47_75 sp47_75 202000.000000
Rwpos47_76 in47_76 sp47_76 78000.000000
Rwpos47_77 in47_77 sp47_77 78000.000000
Rwpos47_78 in47_78 sp47_78 78000.000000
Rwpos47_79 in47_79 sp47_79 78000.000000
Rwpos47_80 in47_80 sp47_80 202000.000000
Rwpos47_81 in47_81 sp47_81 202000.000000
Rwpos47_82 in47_82 sp47_82 78000.000000
Rwpos47_83 in47_83 sp47_83 78000.000000
Rwpos47_84 in47_84 sp47_84 78000.000000
Rwpos48_1 in48_1 sp48_1 78000.000000
Rwpos48_2 in48_2 sp48_2 202000.000000
Rwpos48_3 in48_3 sp48_3 78000.000000
Rwpos48_4 in48_4 sp48_4 78000.000000
Rwpos48_5 in48_5 sp48_5 202000.000000
Rwpos48_6 in48_6 sp48_6 202000.000000
Rwpos48_7 in48_7 sp48_7 202000.000000
Rwpos48_8 in48_8 sp48_8 202000.000000
Rwpos48_9 in48_9 sp48_9 78000.000000
Rwpos48_10 in48_10 sp48_10 78000.000000
Rwpos48_11 in48_11 sp48_11 78000.000000
Rwpos48_12 in48_12 sp48_12 78000.000000
Rwpos48_13 in48_13 sp48_13 78000.000000
Rwpos48_14 in48_14 sp48_14 202000.000000
Rwpos48_15 in48_15 sp48_15 202000.000000
Rwpos48_16 in48_16 sp48_16 202000.000000
Rwpos48_17 in48_17 sp48_17 78000.000000
Rwpos48_18 in48_18 sp48_18 202000.000000
Rwpos48_19 in48_19 sp48_19 78000.000000
Rwpos48_20 in48_20 sp48_20 202000.000000
Rwpos48_21 in48_21 sp48_21 202000.000000
Rwpos48_22 in48_22 sp48_22 78000.000000
Rwpos48_23 in48_23 sp48_23 78000.000000
Rwpos48_24 in48_24 sp48_24 202000.000000
Rwpos48_25 in48_25 sp48_25 78000.000000
Rwpos48_26 in48_26 sp48_26 78000.000000
Rwpos48_27 in48_27 sp48_27 78000.000000
Rwpos48_28 in48_28 sp48_28 78000.000000
Rwpos48_29 in48_29 sp48_29 202000.000000
Rwpos48_30 in48_30 sp48_30 78000.000000
Rwpos48_31 in48_31 sp48_31 78000.000000
Rwpos48_32 in48_32 sp48_32 78000.000000
Rwpos48_33 in48_33 sp48_33 78000.000000
Rwpos48_34 in48_34 sp48_34 78000.000000
Rwpos48_35 in48_35 sp48_35 78000.000000
Rwpos48_36 in48_36 sp48_36 202000.000000
Rwpos48_37 in48_37 sp48_37 78000.000000
Rwpos48_38 in48_38 sp48_38 202000.000000
Rwpos48_39 in48_39 sp48_39 78000.000000
Rwpos48_40 in48_40 sp48_40 78000.000000
Rwpos48_41 in48_41 sp48_41 78000.000000
Rwpos48_42 in48_42 sp48_42 202000.000000
Rwpos48_43 in48_43 sp48_43 202000.000000
Rwpos48_44 in48_44 sp48_44 202000.000000
Rwpos48_45 in48_45 sp48_45 202000.000000
Rwpos48_46 in48_46 sp48_46 78000.000000
Rwpos48_47 in48_47 sp48_47 202000.000000
Rwpos48_48 in48_48 sp48_48 78000.000000
Rwpos48_49 in48_49 sp48_49 202000.000000
Rwpos48_50 in48_50 sp48_50 202000.000000
Rwpos48_51 in48_51 sp48_51 78000.000000
Rwpos48_52 in48_52 sp48_52 202000.000000
Rwpos48_53 in48_53 sp48_53 202000.000000
Rwpos48_54 in48_54 sp48_54 202000.000000
Rwpos48_55 in48_55 sp48_55 78000.000000
Rwpos48_56 in48_56 sp48_56 78000.000000
Rwpos48_57 in48_57 sp48_57 78000.000000
Rwpos48_58 in48_58 sp48_58 78000.000000
Rwpos48_59 in48_59 sp48_59 78000.000000
Rwpos48_60 in48_60 sp48_60 202000.000000
Rwpos48_61 in48_61 sp48_61 78000.000000
Rwpos48_62 in48_62 sp48_62 78000.000000
Rwpos48_63 in48_63 sp48_63 202000.000000
Rwpos48_64 in48_64 sp48_64 202000.000000
Rwpos48_65 in48_65 sp48_65 202000.000000
Rwpos48_66 in48_66 sp48_66 78000.000000
Rwpos48_67 in48_67 sp48_67 78000.000000
Rwpos48_68 in48_68 sp48_68 202000.000000
Rwpos48_69 in48_69 sp48_69 78000.000000
Rwpos48_70 in48_70 sp48_70 78000.000000
Rwpos48_71 in48_71 sp48_71 78000.000000
Rwpos48_72 in48_72 sp48_72 78000.000000
Rwpos48_73 in48_73 sp48_73 78000.000000
Rwpos48_74 in48_74 sp48_74 78000.000000
Rwpos48_75 in48_75 sp48_75 78000.000000
Rwpos48_76 in48_76 sp48_76 202000.000000
Rwpos48_77 in48_77 sp48_77 78000.000000
Rwpos48_78 in48_78 sp48_78 202000.000000
Rwpos48_79 in48_79 sp48_79 78000.000000
Rwpos48_80 in48_80 sp48_80 78000.000000
Rwpos48_81 in48_81 sp48_81 202000.000000
Rwpos48_82 in48_82 sp48_82 202000.000000
Rwpos48_83 in48_83 sp48_83 202000.000000
Rwpos48_84 in48_84 sp48_84 202000.000000
Rwpos49_1 in49_1 sp49_1 78000.000000
Rwpos49_2 in49_2 sp49_2 202000.000000
Rwpos49_3 in49_3 sp49_3 78000.000000
Rwpos49_4 in49_4 sp49_4 202000.000000
Rwpos49_5 in49_5 sp49_5 78000.000000
Rwpos49_6 in49_6 sp49_6 202000.000000
Rwpos49_7 in49_7 sp49_7 202000.000000
Rwpos49_8 in49_8 sp49_8 78000.000000
Rwpos49_9 in49_9 sp49_9 78000.000000
Rwpos49_10 in49_10 sp49_10 78000.000000
Rwpos49_11 in49_11 sp49_11 202000.000000
Rwpos49_12 in49_12 sp49_12 78000.000000
Rwpos49_13 in49_13 sp49_13 78000.000000
Rwpos49_14 in49_14 sp49_14 78000.000000
Rwpos49_15 in49_15 sp49_15 78000.000000
Rwpos49_16 in49_16 sp49_16 78000.000000
Rwpos49_17 in49_17 sp49_17 202000.000000
Rwpos49_18 in49_18 sp49_18 78000.000000
Rwpos49_19 in49_19 sp49_19 78000.000000
Rwpos49_20 in49_20 sp49_20 78000.000000
Rwpos49_21 in49_21 sp49_21 78000.000000
Rwpos49_22 in49_22 sp49_22 78000.000000
Rwpos49_23 in49_23 sp49_23 78000.000000
Rwpos49_24 in49_24 sp49_24 202000.000000
Rwpos49_25 in49_25 sp49_25 202000.000000
Rwpos49_26 in49_26 sp49_26 202000.000000
Rwpos49_27 in49_27 sp49_27 78000.000000
Rwpos49_28 in49_28 sp49_28 78000.000000
Rwpos49_29 in49_29 sp49_29 78000.000000
Rwpos49_30 in49_30 sp49_30 202000.000000
Rwpos49_31 in49_31 sp49_31 78000.000000
Rwpos49_32 in49_32 sp49_32 202000.000000
Rwpos49_33 in49_33 sp49_33 78000.000000
Rwpos49_34 in49_34 sp49_34 202000.000000
Rwpos49_35 in49_35 sp49_35 78000.000000
Rwpos49_36 in49_36 sp49_36 78000.000000
Rwpos49_37 in49_37 sp49_37 202000.000000
Rwpos49_38 in49_38 sp49_38 78000.000000
Rwpos49_39 in49_39 sp49_39 78000.000000
Rwpos49_40 in49_40 sp49_40 78000.000000
Rwpos49_41 in49_41 sp49_41 78000.000000
Rwpos49_42 in49_42 sp49_42 202000.000000
Rwpos49_43 in49_43 sp49_43 78000.000000
Rwpos49_44 in49_44 sp49_44 202000.000000
Rwpos49_45 in49_45 sp49_45 78000.000000
Rwpos49_46 in49_46 sp49_46 202000.000000
Rwpos49_47 in49_47 sp49_47 202000.000000
Rwpos49_48 in49_48 sp49_48 202000.000000
Rwpos49_49 in49_49 sp49_49 78000.000000
Rwpos49_50 in49_50 sp49_50 202000.000000
Rwpos49_51 in49_51 sp49_51 202000.000000
Rwpos49_52 in49_52 sp49_52 78000.000000
Rwpos49_53 in49_53 sp49_53 202000.000000
Rwpos49_54 in49_54 sp49_54 78000.000000
Rwpos49_55 in49_55 sp49_55 202000.000000
Rwpos49_56 in49_56 sp49_56 202000.000000
Rwpos49_57 in49_57 sp49_57 78000.000000
Rwpos49_58 in49_58 sp49_58 78000.000000
Rwpos49_59 in49_59 sp49_59 78000.000000
Rwpos49_60 in49_60 sp49_60 202000.000000
Rwpos49_61 in49_61 sp49_61 78000.000000
Rwpos49_62 in49_62 sp49_62 202000.000000
Rwpos49_63 in49_63 sp49_63 202000.000000
Rwpos49_64 in49_64 sp49_64 202000.000000
Rwpos49_65 in49_65 sp49_65 202000.000000
Rwpos49_66 in49_66 sp49_66 78000.000000
Rwpos49_67 in49_67 sp49_67 78000.000000
Rwpos49_68 in49_68 sp49_68 202000.000000
Rwpos49_69 in49_69 sp49_69 202000.000000
Rwpos49_70 in49_70 sp49_70 78000.000000
Rwpos49_71 in49_71 sp49_71 202000.000000
Rwpos49_72 in49_72 sp49_72 78000.000000
Rwpos49_73 in49_73 sp49_73 78000.000000
Rwpos49_74 in49_74 sp49_74 78000.000000
Rwpos49_75 in49_75 sp49_75 78000.000000
Rwpos49_76 in49_76 sp49_76 78000.000000
Rwpos49_77 in49_77 sp49_77 202000.000000
Rwpos49_78 in49_78 sp49_78 202000.000000
Rwpos49_79 in49_79 sp49_79 202000.000000
Rwpos49_80 in49_80 sp49_80 202000.000000
Rwpos49_81 in49_81 sp49_81 202000.000000
Rwpos49_82 in49_82 sp49_82 78000.000000
Rwpos49_83 in49_83 sp49_83 78000.000000
Rwpos49_84 in49_84 sp49_84 202000.000000
Rwpos50_1 in50_1 sp50_1 78000.000000
Rwpos50_2 in50_2 sp50_2 78000.000000
Rwpos50_3 in50_3 sp50_3 78000.000000
Rwpos50_4 in50_4 sp50_4 202000.000000
Rwpos50_5 in50_5 sp50_5 78000.000000
Rwpos50_6 in50_6 sp50_6 78000.000000
Rwpos50_7 in50_7 sp50_7 202000.000000
Rwpos50_8 in50_8 sp50_8 78000.000000
Rwpos50_9 in50_9 sp50_9 78000.000000
Rwpos50_10 in50_10 sp50_10 78000.000000
Rwpos50_11 in50_11 sp50_11 78000.000000
Rwpos50_12 in50_12 sp50_12 202000.000000
Rwpos50_13 in50_13 sp50_13 78000.000000
Rwpos50_14 in50_14 sp50_14 78000.000000
Rwpos50_15 in50_15 sp50_15 78000.000000
Rwpos50_16 in50_16 sp50_16 202000.000000
Rwpos50_17 in50_17 sp50_17 78000.000000
Rwpos50_18 in50_18 sp50_18 202000.000000
Rwpos50_19 in50_19 sp50_19 202000.000000
Rwpos50_20 in50_20 sp50_20 78000.000000
Rwpos50_21 in50_21 sp50_21 78000.000000
Rwpos50_22 in50_22 sp50_22 78000.000000
Rwpos50_23 in50_23 sp50_23 202000.000000
Rwpos50_24 in50_24 sp50_24 78000.000000
Rwpos50_25 in50_25 sp50_25 78000.000000
Rwpos50_26 in50_26 sp50_26 78000.000000
Rwpos50_27 in50_27 sp50_27 78000.000000
Rwpos50_28 in50_28 sp50_28 202000.000000
Rwpos50_29 in50_29 sp50_29 202000.000000
Rwpos50_30 in50_30 sp50_30 78000.000000
Rwpos50_31 in50_31 sp50_31 78000.000000
Rwpos50_32 in50_32 sp50_32 78000.000000
Rwpos50_33 in50_33 sp50_33 78000.000000
Rwpos50_34 in50_34 sp50_34 78000.000000
Rwpos50_35 in50_35 sp50_35 78000.000000
Rwpos50_36 in50_36 sp50_36 78000.000000
Rwpos50_37 in50_37 sp50_37 202000.000000
Rwpos50_38 in50_38 sp50_38 202000.000000
Rwpos50_39 in50_39 sp50_39 202000.000000
Rwpos50_40 in50_40 sp50_40 202000.000000
Rwpos50_41 in50_41 sp50_41 78000.000000
Rwpos50_42 in50_42 sp50_42 202000.000000
Rwpos50_43 in50_43 sp50_43 202000.000000
Rwpos50_44 in50_44 sp50_44 202000.000000
Rwpos50_45 in50_45 sp50_45 78000.000000
Rwpos50_46 in50_46 sp50_46 78000.000000
Rwpos50_47 in50_47 sp50_47 202000.000000
Rwpos50_48 in50_48 sp50_48 202000.000000
Rwpos50_49 in50_49 sp50_49 78000.000000
Rwpos50_50 in50_50 sp50_50 78000.000000
Rwpos50_51 in50_51 sp50_51 202000.000000
Rwpos50_52 in50_52 sp50_52 78000.000000
Rwpos50_53 in50_53 sp50_53 78000.000000
Rwpos50_54 in50_54 sp50_54 202000.000000
Rwpos50_55 in50_55 sp50_55 78000.000000
Rwpos50_56 in50_56 sp50_56 202000.000000
Rwpos50_57 in50_57 sp50_57 78000.000000
Rwpos50_58 in50_58 sp50_58 78000.000000
Rwpos50_59 in50_59 sp50_59 78000.000000
Rwpos50_60 in50_60 sp50_60 202000.000000
Rwpos50_61 in50_61 sp50_61 78000.000000
Rwpos50_62 in50_62 sp50_62 202000.000000
Rwpos50_63 in50_63 sp50_63 78000.000000
Rwpos50_64 in50_64 sp50_64 78000.000000
Rwpos50_65 in50_65 sp50_65 202000.000000
Rwpos50_66 in50_66 sp50_66 202000.000000
Rwpos50_67 in50_67 sp50_67 78000.000000
Rwpos50_68 in50_68 sp50_68 202000.000000
Rwpos50_69 in50_69 sp50_69 202000.000000
Rwpos50_70 in50_70 sp50_70 78000.000000
Rwpos50_71 in50_71 sp50_71 202000.000000
Rwpos50_72 in50_72 sp50_72 78000.000000
Rwpos50_73 in50_73 sp50_73 78000.000000
Rwpos50_74 in50_74 sp50_74 78000.000000
Rwpos50_75 in50_75 sp50_75 78000.000000
Rwpos50_76 in50_76 sp50_76 78000.000000
Rwpos50_77 in50_77 sp50_77 202000.000000
Rwpos50_78 in50_78 sp50_78 78000.000000
Rwpos50_79 in50_79 sp50_79 202000.000000
Rwpos50_80 in50_80 sp50_80 78000.000000
Rwpos50_81 in50_81 sp50_81 202000.000000
Rwpos50_82 in50_82 sp50_82 78000.000000
Rwpos50_83 in50_83 sp50_83 78000.000000
Rwpos50_84 in50_84 sp50_84 78000.000000
Rwpos51_1 in51_1 sp51_1 78000.000000
Rwpos51_2 in51_2 sp51_2 78000.000000
Rwpos51_3 in51_3 sp51_3 202000.000000
Rwpos51_4 in51_4 sp51_4 78000.000000
Rwpos51_5 in51_5 sp51_5 202000.000000
Rwpos51_6 in51_6 sp51_6 78000.000000
Rwpos51_7 in51_7 sp51_7 202000.000000
Rwpos51_8 in51_8 sp51_8 202000.000000
Rwpos51_9 in51_9 sp51_9 202000.000000
Rwpos51_10 in51_10 sp51_10 78000.000000
Rwpos51_11 in51_11 sp51_11 202000.000000
Rwpos51_12 in51_12 sp51_12 78000.000000
Rwpos51_13 in51_13 sp51_13 202000.000000
Rwpos51_14 in51_14 sp51_14 78000.000000
Rwpos51_15 in51_15 sp51_15 78000.000000
Rwpos51_16 in51_16 sp51_16 78000.000000
Rwpos51_17 in51_17 sp51_17 78000.000000
Rwpos51_18 in51_18 sp51_18 202000.000000
Rwpos51_19 in51_19 sp51_19 78000.000000
Rwpos51_20 in51_20 sp51_20 202000.000000
Rwpos51_21 in51_21 sp51_21 78000.000000
Rwpos51_22 in51_22 sp51_22 78000.000000
Rwpos51_23 in51_23 sp51_23 202000.000000
Rwpos51_24 in51_24 sp51_24 78000.000000
Rwpos51_25 in51_25 sp51_25 202000.000000
Rwpos51_26 in51_26 sp51_26 78000.000000
Rwpos51_27 in51_27 sp51_27 202000.000000
Rwpos51_28 in51_28 sp51_28 78000.000000
Rwpos51_29 in51_29 sp51_29 202000.000000
Rwpos51_30 in51_30 sp51_30 78000.000000
Rwpos51_31 in51_31 sp51_31 78000.000000
Rwpos51_32 in51_32 sp51_32 202000.000000
Rwpos51_33 in51_33 sp51_33 78000.000000
Rwpos51_34 in51_34 sp51_34 202000.000000
Rwpos51_35 in51_35 sp51_35 202000.000000
Rwpos51_36 in51_36 sp51_36 202000.000000
Rwpos51_37 in51_37 sp51_37 202000.000000
Rwpos51_38 in51_38 sp51_38 78000.000000
Rwpos51_39 in51_39 sp51_39 78000.000000
Rwpos51_40 in51_40 sp51_40 78000.000000
Rwpos51_41 in51_41 sp51_41 202000.000000
Rwpos51_42 in51_42 sp51_42 202000.000000
Rwpos51_43 in51_43 sp51_43 202000.000000
Rwpos51_44 in51_44 sp51_44 78000.000000
Rwpos51_45 in51_45 sp51_45 78000.000000
Rwpos51_46 in51_46 sp51_46 202000.000000
Rwpos51_47 in51_47 sp51_47 78000.000000
Rwpos51_48 in51_48 sp51_48 202000.000000
Rwpos51_49 in51_49 sp51_49 202000.000000
Rwpos51_50 in51_50 sp51_50 78000.000000
Rwpos51_51 in51_51 sp51_51 78000.000000
Rwpos51_52 in51_52 sp51_52 78000.000000
Rwpos51_53 in51_53 sp51_53 78000.000000
Rwpos51_54 in51_54 sp51_54 78000.000000
Rwpos51_55 in51_55 sp51_55 202000.000000
Rwpos51_56 in51_56 sp51_56 202000.000000
Rwpos51_57 in51_57 sp51_57 78000.000000
Rwpos51_58 in51_58 sp51_58 202000.000000
Rwpos51_59 in51_59 sp51_59 202000.000000
Rwpos51_60 in51_60 sp51_60 202000.000000
Rwpos51_61 in51_61 sp51_61 78000.000000
Rwpos51_62 in51_62 sp51_62 202000.000000
Rwpos51_63 in51_63 sp51_63 78000.000000
Rwpos51_64 in51_64 sp51_64 202000.000000
Rwpos51_65 in51_65 sp51_65 202000.000000
Rwpos51_66 in51_66 sp51_66 202000.000000
Rwpos51_67 in51_67 sp51_67 78000.000000
Rwpos51_68 in51_68 sp51_68 78000.000000
Rwpos51_69 in51_69 sp51_69 202000.000000
Rwpos51_70 in51_70 sp51_70 78000.000000
Rwpos51_71 in51_71 sp51_71 202000.000000
Rwpos51_72 in51_72 sp51_72 78000.000000
Rwpos51_73 in51_73 sp51_73 78000.000000
Rwpos51_74 in51_74 sp51_74 78000.000000
Rwpos51_75 in51_75 sp51_75 202000.000000
Rwpos51_76 in51_76 sp51_76 202000.000000
Rwpos51_77 in51_77 sp51_77 78000.000000
Rwpos51_78 in51_78 sp51_78 78000.000000
Rwpos51_79 in51_79 sp51_79 202000.000000
Rwpos51_80 in51_80 sp51_80 202000.000000
Rwpos51_81 in51_81 sp51_81 202000.000000
Rwpos51_82 in51_82 sp51_82 78000.000000
Rwpos51_83 in51_83 sp51_83 78000.000000
Rwpos51_84 in51_84 sp51_84 78000.000000
Rwpos52_1 in52_1 sp52_1 202000.000000
Rwpos52_2 in52_2 sp52_2 202000.000000
Rwpos52_3 in52_3 sp52_3 78000.000000
Rwpos52_4 in52_4 sp52_4 78000.000000
Rwpos52_5 in52_5 sp52_5 202000.000000
Rwpos52_6 in52_6 sp52_6 202000.000000
Rwpos52_7 in52_7 sp52_7 202000.000000
Rwpos52_8 in52_8 sp52_8 78000.000000
Rwpos52_9 in52_9 sp52_9 78000.000000
Rwpos52_10 in52_10 sp52_10 202000.000000
Rwpos52_11 in52_11 sp52_11 78000.000000
Rwpos52_12 in52_12 sp52_12 78000.000000
Rwpos52_13 in52_13 sp52_13 78000.000000
Rwpos52_14 in52_14 sp52_14 202000.000000
Rwpos52_15 in52_15 sp52_15 78000.000000
Rwpos52_16 in52_16 sp52_16 78000.000000
Rwpos52_17 in52_17 sp52_17 78000.000000
Rwpos52_18 in52_18 sp52_18 202000.000000
Rwpos52_19 in52_19 sp52_19 78000.000000
Rwpos52_20 in52_20 sp52_20 78000.000000
Rwpos52_21 in52_21 sp52_21 202000.000000
Rwpos52_22 in52_22 sp52_22 78000.000000
Rwpos52_23 in52_23 sp52_23 78000.000000
Rwpos52_24 in52_24 sp52_24 202000.000000
Rwpos52_25 in52_25 sp52_25 78000.000000
Rwpos52_26 in52_26 sp52_26 78000.000000
Rwpos52_27 in52_27 sp52_27 202000.000000
Rwpos52_28 in52_28 sp52_28 78000.000000
Rwpos52_29 in52_29 sp52_29 202000.000000
Rwpos52_30 in52_30 sp52_30 78000.000000
Rwpos52_31 in52_31 sp52_31 78000.000000
Rwpos52_32 in52_32 sp52_32 202000.000000
Rwpos52_33 in52_33 sp52_33 78000.000000
Rwpos52_34 in52_34 sp52_34 202000.000000
Rwpos52_35 in52_35 sp52_35 78000.000000
Rwpos52_36 in52_36 sp52_36 202000.000000
Rwpos52_37 in52_37 sp52_37 202000.000000
Rwpos52_38 in52_38 sp52_38 78000.000000
Rwpos52_39 in52_39 sp52_39 78000.000000
Rwpos52_40 in52_40 sp52_40 78000.000000
Rwpos52_41 in52_41 sp52_41 78000.000000
Rwpos52_42 in52_42 sp52_42 202000.000000
Rwpos52_43 in52_43 sp52_43 78000.000000
Rwpos52_44 in52_44 sp52_44 202000.000000
Rwpos52_45 in52_45 sp52_45 78000.000000
Rwpos52_46 in52_46 sp52_46 202000.000000
Rwpos52_47 in52_47 sp52_47 202000.000000
Rwpos52_48 in52_48 sp52_48 202000.000000
Rwpos52_49 in52_49 sp52_49 78000.000000
Rwpos52_50 in52_50 sp52_50 202000.000000
Rwpos52_51 in52_51 sp52_51 78000.000000
Rwpos52_52 in52_52 sp52_52 202000.000000
Rwpos52_53 in52_53 sp52_53 78000.000000
Rwpos52_54 in52_54 sp52_54 202000.000000
Rwpos52_55 in52_55 sp52_55 202000.000000
Rwpos52_56 in52_56 sp52_56 78000.000000
Rwpos52_57 in52_57 sp52_57 78000.000000
Rwpos52_58 in52_58 sp52_58 78000.000000
Rwpos52_59 in52_59 sp52_59 78000.000000
Rwpos52_60 in52_60 sp52_60 202000.000000
Rwpos52_61 in52_61 sp52_61 78000.000000
Rwpos52_62 in52_62 sp52_62 202000.000000
Rwpos52_63 in52_63 sp52_63 78000.000000
Rwpos52_64 in52_64 sp52_64 78000.000000
Rwpos52_65 in52_65 sp52_65 202000.000000
Rwpos52_66 in52_66 sp52_66 202000.000000
Rwpos52_67 in52_67 sp52_67 202000.000000
Rwpos52_68 in52_68 sp52_68 202000.000000
Rwpos52_69 in52_69 sp52_69 202000.000000
Rwpos52_70 in52_70 sp52_70 78000.000000
Rwpos52_71 in52_71 sp52_71 202000.000000
Rwpos52_72 in52_72 sp52_72 78000.000000
Rwpos52_73 in52_73 sp52_73 202000.000000
Rwpos52_74 in52_74 sp52_74 78000.000000
Rwpos52_75 in52_75 sp52_75 78000.000000
Rwpos52_76 in52_76 sp52_76 78000.000000
Rwpos52_77 in52_77 sp52_77 202000.000000
Rwpos52_78 in52_78 sp52_78 78000.000000
Rwpos52_79 in52_79 sp52_79 202000.000000
Rwpos52_80 in52_80 sp52_80 78000.000000
Rwpos52_81 in52_81 sp52_81 202000.000000
Rwpos52_82 in52_82 sp52_82 202000.000000
Rwpos52_83 in52_83 sp52_83 78000.000000
Rwpos52_84 in52_84 sp52_84 78000.000000
Rwpos53_1 in53_1 sp53_1 78000.000000
Rwpos53_2 in53_2 sp53_2 202000.000000
Rwpos53_3 in53_3 sp53_3 78000.000000
Rwpos53_4 in53_4 sp53_4 202000.000000
Rwpos53_5 in53_5 sp53_5 202000.000000
Rwpos53_6 in53_6 sp53_6 78000.000000
Rwpos53_7 in53_7 sp53_7 78000.000000
Rwpos53_8 in53_8 sp53_8 202000.000000
Rwpos53_9 in53_9 sp53_9 202000.000000
Rwpos53_10 in53_10 sp53_10 78000.000000
Rwpos53_11 in53_11 sp53_11 202000.000000
Rwpos53_12 in53_12 sp53_12 202000.000000
Rwpos53_13 in53_13 sp53_13 78000.000000
Rwpos53_14 in53_14 sp53_14 202000.000000
Rwpos53_15 in53_15 sp53_15 78000.000000
Rwpos53_16 in53_16 sp53_16 202000.000000
Rwpos53_17 in53_17 sp53_17 78000.000000
Rwpos53_18 in53_18 sp53_18 78000.000000
Rwpos53_19 in53_19 sp53_19 78000.000000
Rwpos53_20 in53_20 sp53_20 78000.000000
Rwpos53_21 in53_21 sp53_21 78000.000000
Rwpos53_22 in53_22 sp53_22 202000.000000
Rwpos53_23 in53_23 sp53_23 78000.000000
Rwpos53_24 in53_24 sp53_24 78000.000000
Rwpos53_25 in53_25 sp53_25 202000.000000
Rwpos53_26 in53_26 sp53_26 78000.000000
Rwpos53_27 in53_27 sp53_27 202000.000000
Rwpos53_28 in53_28 sp53_28 78000.000000
Rwpos53_29 in53_29 sp53_29 78000.000000
Rwpos53_30 in53_30 sp53_30 202000.000000
Rwpos53_31 in53_31 sp53_31 202000.000000
Rwpos53_32 in53_32 sp53_32 78000.000000
Rwpos53_33 in53_33 sp53_33 78000.000000
Rwpos53_34 in53_34 sp53_34 202000.000000
Rwpos53_35 in53_35 sp53_35 202000.000000
Rwpos53_36 in53_36 sp53_36 202000.000000
Rwpos53_37 in53_37 sp53_37 78000.000000
Rwpos53_38 in53_38 sp53_38 78000.000000
Rwpos53_39 in53_39 sp53_39 78000.000000
Rwpos53_40 in53_40 sp53_40 78000.000000
Rwpos53_41 in53_41 sp53_41 202000.000000
Rwpos53_42 in53_42 sp53_42 78000.000000
Rwpos53_43 in53_43 sp53_43 78000.000000
Rwpos53_44 in53_44 sp53_44 202000.000000
Rwpos53_45 in53_45 sp53_45 78000.000000
Rwpos53_46 in53_46 sp53_46 202000.000000
Rwpos53_47 in53_47 sp53_47 202000.000000
Rwpos53_48 in53_48 sp53_48 202000.000000
Rwpos53_49 in53_49 sp53_49 202000.000000
Rwpos53_50 in53_50 sp53_50 78000.000000
Rwpos53_51 in53_51 sp53_51 202000.000000
Rwpos53_52 in53_52 sp53_52 202000.000000
Rwpos53_53 in53_53 sp53_53 202000.000000
Rwpos53_54 in53_54 sp53_54 78000.000000
Rwpos53_55 in53_55 sp53_55 202000.000000
Rwpos53_56 in53_56 sp53_56 78000.000000
Rwpos53_57 in53_57 sp53_57 202000.000000
Rwpos53_58 in53_58 sp53_58 78000.000000
Rwpos53_59 in53_59 sp53_59 78000.000000
Rwpos53_60 in53_60 sp53_60 202000.000000
Rwpos53_61 in53_61 sp53_61 202000.000000
Rwpos53_62 in53_62 sp53_62 78000.000000
Rwpos53_63 in53_63 sp53_63 202000.000000
Rwpos53_64 in53_64 sp53_64 202000.000000
Rwpos53_65 in53_65 sp53_65 78000.000000
Rwpos53_66 in53_66 sp53_66 78000.000000
Rwpos53_67 in53_67 sp53_67 202000.000000
Rwpos53_68 in53_68 sp53_68 78000.000000
Rwpos53_69 in53_69 sp53_69 202000.000000
Rwpos53_70 in53_70 sp53_70 202000.000000
Rwpos53_71 in53_71 sp53_71 78000.000000
Rwpos53_72 in53_72 sp53_72 202000.000000
Rwpos53_73 in53_73 sp53_73 202000.000000
Rwpos53_74 in53_74 sp53_74 202000.000000
Rwpos53_75 in53_75 sp53_75 202000.000000
Rwpos53_76 in53_76 sp53_76 202000.000000
Rwpos53_77 in53_77 sp53_77 78000.000000
Rwpos53_78 in53_78 sp53_78 78000.000000
Rwpos53_79 in53_79 sp53_79 78000.000000
Rwpos53_80 in53_80 sp53_80 78000.000000
Rwpos53_81 in53_81 sp53_81 78000.000000
Rwpos53_82 in53_82 sp53_82 202000.000000
Rwpos53_83 in53_83 sp53_83 78000.000000
Rwpos53_84 in53_84 sp53_84 78000.000000
Rwpos54_1 in54_1 sp54_1 202000.000000
Rwpos54_2 in54_2 sp54_2 78000.000000
Rwpos54_3 in54_3 sp54_3 78000.000000
Rwpos54_4 in54_4 sp54_4 202000.000000
Rwpos54_5 in54_5 sp54_5 202000.000000
Rwpos54_6 in54_6 sp54_6 78000.000000
Rwpos54_7 in54_7 sp54_7 78000.000000
Rwpos54_8 in54_8 sp54_8 78000.000000
Rwpos54_9 in54_9 sp54_9 78000.000000
Rwpos54_10 in54_10 sp54_10 78000.000000
Rwpos54_11 in54_11 sp54_11 78000.000000
Rwpos54_12 in54_12 sp54_12 202000.000000
Rwpos54_13 in54_13 sp54_13 202000.000000
Rwpos54_14 in54_14 sp54_14 78000.000000
Rwpos54_15 in54_15 sp54_15 202000.000000
Rwpos54_16 in54_16 sp54_16 202000.000000
Rwpos54_17 in54_17 sp54_17 78000.000000
Rwpos54_18 in54_18 sp54_18 202000.000000
Rwpos54_19 in54_19 sp54_19 202000.000000
Rwpos54_20 in54_20 sp54_20 202000.000000
Rwpos54_21 in54_21 sp54_21 78000.000000
Rwpos54_22 in54_22 sp54_22 202000.000000
Rwpos54_23 in54_23 sp54_23 78000.000000
Rwpos54_24 in54_24 sp54_24 202000.000000
Rwpos54_25 in54_25 sp54_25 78000.000000
Rwpos54_26 in54_26 sp54_26 202000.000000
Rwpos54_27 in54_27 sp54_27 202000.000000
Rwpos54_28 in54_28 sp54_28 202000.000000
Rwpos54_29 in54_29 sp54_29 78000.000000
Rwpos54_30 in54_30 sp54_30 78000.000000
Rwpos54_31 in54_31 sp54_31 202000.000000
Rwpos54_32 in54_32 sp54_32 202000.000000
Rwpos54_33 in54_33 sp54_33 78000.000000
Rwpos54_34 in54_34 sp54_34 78000.000000
Rwpos54_35 in54_35 sp54_35 78000.000000
Rwpos54_36 in54_36 sp54_36 78000.000000
Rwpos54_37 in54_37 sp54_37 78000.000000
Rwpos54_38 in54_38 sp54_38 202000.000000
Rwpos54_39 in54_39 sp54_39 202000.000000
Rwpos54_40 in54_40 sp54_40 202000.000000
Rwpos54_41 in54_41 sp54_41 202000.000000
Rwpos54_42 in54_42 sp54_42 78000.000000
Rwpos54_43 in54_43 sp54_43 78000.000000
Rwpos54_44 in54_44 sp54_44 78000.000000
Rwpos54_45 in54_45 sp54_45 202000.000000
Rwpos54_46 in54_46 sp54_46 202000.000000
Rwpos54_47 in54_47 sp54_47 78000.000000
Rwpos54_48 in54_48 sp54_48 202000.000000
Rwpos54_49 in54_49 sp54_49 78000.000000
Rwpos54_50 in54_50 sp54_50 78000.000000
Rwpos54_51 in54_51 sp54_51 202000.000000
Rwpos54_52 in54_52 sp54_52 78000.000000
Rwpos54_53 in54_53 sp54_53 202000.000000
Rwpos54_54 in54_54 sp54_54 202000.000000
Rwpos54_55 in54_55 sp54_55 202000.000000
Rwpos54_56 in54_56 sp54_56 202000.000000
Rwpos54_57 in54_57 sp54_57 78000.000000
Rwpos54_58 in54_58 sp54_58 78000.000000
Rwpos54_59 in54_59 sp54_59 78000.000000
Rwpos54_60 in54_60 sp54_60 78000.000000
Rwpos54_61 in54_61 sp54_61 78000.000000
Rwpos54_62 in54_62 sp54_62 202000.000000
Rwpos54_63 in54_63 sp54_63 78000.000000
Rwpos54_64 in54_64 sp54_64 202000.000000
Rwpos54_65 in54_65 sp54_65 78000.000000
Rwpos54_66 in54_66 sp54_66 202000.000000
Rwpos54_67 in54_67 sp54_67 202000.000000
Rwpos54_68 in54_68 sp54_68 78000.000000
Rwpos54_69 in54_69 sp54_69 202000.000000
Rwpos54_70 in54_70 sp54_70 202000.000000
Rwpos54_71 in54_71 sp54_71 78000.000000
Rwpos54_72 in54_72 sp54_72 78000.000000
Rwpos54_73 in54_73 sp54_73 78000.000000
Rwpos54_74 in54_74 sp54_74 78000.000000
Rwpos54_75 in54_75 sp54_75 202000.000000
Rwpos54_76 in54_76 sp54_76 78000.000000
Rwpos54_77 in54_77 sp54_77 78000.000000
Rwpos54_78 in54_78 sp54_78 202000.000000
Rwpos54_79 in54_79 sp54_79 202000.000000
Rwpos54_80 in54_80 sp54_80 202000.000000
Rwpos54_81 in54_81 sp54_81 78000.000000
Rwpos54_82 in54_82 sp54_82 78000.000000
Rwpos54_83 in54_83 sp54_83 78000.000000
Rwpos54_84 in54_84 sp54_84 78000.000000
Rwpos55_1 in55_1 sp55_1 202000.000000
Rwpos55_2 in55_2 sp55_2 202000.000000
Rwpos55_3 in55_3 sp55_3 202000.000000
Rwpos55_4 in55_4 sp55_4 202000.000000
Rwpos55_5 in55_5 sp55_5 202000.000000
Rwpos55_6 in55_6 sp55_6 78000.000000
Rwpos55_7 in55_7 sp55_7 78000.000000
Rwpos55_8 in55_8 sp55_8 202000.000000
Rwpos55_9 in55_9 sp55_9 202000.000000
Rwpos55_10 in55_10 sp55_10 202000.000000
Rwpos55_11 in55_11 sp55_11 78000.000000
Rwpos55_12 in55_12 sp55_12 202000.000000
Rwpos55_13 in55_13 sp55_13 78000.000000
Rwpos55_14 in55_14 sp55_14 78000.000000
Rwpos55_15 in55_15 sp55_15 78000.000000
Rwpos55_16 in55_16 sp55_16 202000.000000
Rwpos55_17 in55_17 sp55_17 78000.000000
Rwpos55_18 in55_18 sp55_18 202000.000000
Rwpos55_19 in55_19 sp55_19 78000.000000
Rwpos55_20 in55_20 sp55_20 202000.000000
Rwpos55_21 in55_21 sp55_21 78000.000000
Rwpos55_22 in55_22 sp55_22 202000.000000
Rwpos55_23 in55_23 sp55_23 78000.000000
Rwpos55_24 in55_24 sp55_24 78000.000000
Rwpos55_25 in55_25 sp55_25 202000.000000
Rwpos55_26 in55_26 sp55_26 202000.000000
Rwpos55_27 in55_27 sp55_27 202000.000000
Rwpos55_28 in55_28 sp55_28 202000.000000
Rwpos55_29 in55_29 sp55_29 78000.000000
Rwpos55_30 in55_30 sp55_30 78000.000000
Rwpos55_31 in55_31 sp55_31 78000.000000
Rwpos55_32 in55_32 sp55_32 78000.000000
Rwpos55_33 in55_33 sp55_33 202000.000000
Rwpos55_34 in55_34 sp55_34 202000.000000
Rwpos55_35 in55_35 sp55_35 78000.000000
Rwpos55_36 in55_36 sp55_36 78000.000000
Rwpos55_37 in55_37 sp55_37 202000.000000
Rwpos55_38 in55_38 sp55_38 78000.000000
Rwpos55_39 in55_39 sp55_39 78000.000000
Rwpos55_40 in55_40 sp55_40 78000.000000
Rwpos55_41 in55_41 sp55_41 78000.000000
Rwpos55_42 in55_42 sp55_42 202000.000000
Rwpos55_43 in55_43 sp55_43 202000.000000
Rwpos55_44 in55_44 sp55_44 78000.000000
Rwpos55_45 in55_45 sp55_45 202000.000000
Rwpos55_46 in55_46 sp55_46 78000.000000
Rwpos55_47 in55_47 sp55_47 78000.000000
Rwpos55_48 in55_48 sp55_48 78000.000000
Rwpos55_49 in55_49 sp55_49 202000.000000
Rwpos55_50 in55_50 sp55_50 202000.000000
Rwpos55_51 in55_51 sp55_51 78000.000000
Rwpos55_52 in55_52 sp55_52 202000.000000
Rwpos55_53 in55_53 sp55_53 78000.000000
Rwpos55_54 in55_54 sp55_54 202000.000000
Rwpos55_55 in55_55 sp55_55 202000.000000
Rwpos55_56 in55_56 sp55_56 78000.000000
Rwpos55_57 in55_57 sp55_57 78000.000000
Rwpos55_58 in55_58 sp55_58 78000.000000
Rwpos55_59 in55_59 sp55_59 78000.000000
Rwpos55_60 in55_60 sp55_60 78000.000000
Rwpos55_61 in55_61 sp55_61 202000.000000
Rwpos55_62 in55_62 sp55_62 78000.000000
Rwpos55_63 in55_63 sp55_63 78000.000000
Rwpos55_64 in55_64 sp55_64 202000.000000
Rwpos55_65 in55_65 sp55_65 78000.000000
Rwpos55_66 in55_66 sp55_66 78000.000000
Rwpos55_67 in55_67 sp55_67 78000.000000
Rwpos55_68 in55_68 sp55_68 78000.000000
Rwpos55_69 in55_69 sp55_69 202000.000000
Rwpos55_70 in55_70 sp55_70 78000.000000
Rwpos55_71 in55_71 sp55_71 202000.000000
Rwpos55_72 in55_72 sp55_72 78000.000000
Rwpos55_73 in55_73 sp55_73 78000.000000
Rwpos55_74 in55_74 sp55_74 78000.000000
Rwpos55_75 in55_75 sp55_75 78000.000000
Rwpos55_76 in55_76 sp55_76 78000.000000
Rwpos55_77 in55_77 sp55_77 78000.000000
Rwpos55_78 in55_78 sp55_78 202000.000000
Rwpos55_79 in55_79 sp55_79 78000.000000
Rwpos55_80 in55_80 sp55_80 202000.000000
Rwpos55_81 in55_81 sp55_81 78000.000000
Rwpos55_82 in55_82 sp55_82 202000.000000
Rwpos55_83 in55_83 sp55_83 202000.000000
Rwpos55_84 in55_84 sp55_84 202000.000000
Rwpos56_1 in56_1 sp56_1 202000.000000
Rwpos56_2 in56_2 sp56_2 78000.000000
Rwpos56_3 in56_3 sp56_3 202000.000000
Rwpos56_4 in56_4 sp56_4 202000.000000
Rwpos56_5 in56_5 sp56_5 78000.000000
Rwpos56_6 in56_6 sp56_6 78000.000000
Rwpos56_7 in56_7 sp56_7 78000.000000
Rwpos56_8 in56_8 sp56_8 78000.000000
Rwpos56_9 in56_9 sp56_9 78000.000000
Rwpos56_10 in56_10 sp56_10 202000.000000
Rwpos56_11 in56_11 sp56_11 202000.000000
Rwpos56_12 in56_12 sp56_12 202000.000000
Rwpos56_13 in56_13 sp56_13 202000.000000
Rwpos56_14 in56_14 sp56_14 202000.000000
Rwpos56_15 in56_15 sp56_15 202000.000000
Rwpos56_16 in56_16 sp56_16 202000.000000
Rwpos56_17 in56_17 sp56_17 78000.000000
Rwpos56_18 in56_18 sp56_18 78000.000000
Rwpos56_19 in56_19 sp56_19 78000.000000
Rwpos56_20 in56_20 sp56_20 202000.000000
Rwpos56_21 in56_21 sp56_21 78000.000000
Rwpos56_22 in56_22 sp56_22 202000.000000
Rwpos56_23 in56_23 sp56_23 78000.000000
Rwpos56_24 in56_24 sp56_24 202000.000000
Rwpos56_25 in56_25 sp56_25 78000.000000
Rwpos56_26 in56_26 sp56_26 78000.000000
Rwpos56_27 in56_27 sp56_27 202000.000000
Rwpos56_28 in56_28 sp56_28 202000.000000
Rwpos56_29 in56_29 sp56_29 202000.000000
Rwpos56_30 in56_30 sp56_30 78000.000000
Rwpos56_31 in56_31 sp56_31 202000.000000
Rwpos56_32 in56_32 sp56_32 78000.000000
Rwpos56_33 in56_33 sp56_33 202000.000000
Rwpos56_34 in56_34 sp56_34 78000.000000
Rwpos56_35 in56_35 sp56_35 202000.000000
Rwpos56_36 in56_36 sp56_36 78000.000000
Rwpos56_37 in56_37 sp56_37 78000.000000
Rwpos56_38 in56_38 sp56_38 202000.000000
Rwpos56_39 in56_39 sp56_39 202000.000000
Rwpos56_40 in56_40 sp56_40 78000.000000
Rwpos56_41 in56_41 sp56_41 202000.000000
Rwpos56_42 in56_42 sp56_42 78000.000000
Rwpos56_43 in56_43 sp56_43 202000.000000
Rwpos56_44 in56_44 sp56_44 78000.000000
Rwpos56_45 in56_45 sp56_45 202000.000000
Rwpos56_46 in56_46 sp56_46 202000.000000
Rwpos56_47 in56_47 sp56_47 202000.000000
Rwpos56_48 in56_48 sp56_48 78000.000000
Rwpos56_49 in56_49 sp56_49 78000.000000
Rwpos56_50 in56_50 sp56_50 202000.000000
Rwpos56_51 in56_51 sp56_51 78000.000000
Rwpos56_52 in56_52 sp56_52 202000.000000
Rwpos56_53 in56_53 sp56_53 78000.000000
Rwpos56_54 in56_54 sp56_54 78000.000000
Rwpos56_55 in56_55 sp56_55 202000.000000
Rwpos56_56 in56_56 sp56_56 78000.000000
Rwpos56_57 in56_57 sp56_57 202000.000000
Rwpos56_58 in56_58 sp56_58 78000.000000
Rwpos56_59 in56_59 sp56_59 78000.000000
Rwpos56_60 in56_60 sp56_60 78000.000000
Rwpos56_61 in56_61 sp56_61 78000.000000
Rwpos56_62 in56_62 sp56_62 78000.000000
Rwpos56_63 in56_63 sp56_63 78000.000000
Rwpos56_64 in56_64 sp56_64 202000.000000
Rwpos56_65 in56_65 sp56_65 78000.000000
Rwpos56_66 in56_66 sp56_66 78000.000000
Rwpos56_67 in56_67 sp56_67 202000.000000
Rwpos56_68 in56_68 sp56_68 78000.000000
Rwpos56_69 in56_69 sp56_69 78000.000000
Rwpos56_70 in56_70 sp56_70 202000.000000
Rwpos56_71 in56_71 sp56_71 78000.000000
Rwpos56_72 in56_72 sp56_72 202000.000000
Rwpos56_73 in56_73 sp56_73 78000.000000
Rwpos56_74 in56_74 sp56_74 202000.000000
Rwpos56_75 in56_75 sp56_75 202000.000000
Rwpos56_76 in56_76 sp56_76 78000.000000
Rwpos56_77 in56_77 sp56_77 78000.000000
Rwpos56_78 in56_78 sp56_78 202000.000000
Rwpos56_79 in56_79 sp56_79 78000.000000
Rwpos56_80 in56_80 sp56_80 78000.000000
Rwpos56_81 in56_81 sp56_81 78000.000000
Rwpos56_82 in56_82 sp56_82 78000.000000
Rwpos56_83 in56_83 sp56_83 78000.000000
Rwpos56_84 in56_84 sp56_84 202000.000000
Rwpos57_1 in57_1 sp57_1 78000.000000
Rwpos57_2 in57_2 sp57_2 202000.000000
Rwpos57_3 in57_3 sp57_3 78000.000000
Rwpos57_4 in57_4 sp57_4 78000.000000
Rwpos57_5 in57_5 sp57_5 78000.000000
Rwpos57_6 in57_6 sp57_6 202000.000000
Rwpos57_7 in57_7 sp57_7 202000.000000
Rwpos57_8 in57_8 sp57_8 202000.000000
Rwpos57_9 in57_9 sp57_9 78000.000000
Rwpos57_10 in57_10 sp57_10 202000.000000
Rwpos57_11 in57_11 sp57_11 78000.000000
Rwpos57_12 in57_12 sp57_12 78000.000000
Rwpos57_13 in57_13 sp57_13 202000.000000
Rwpos57_14 in57_14 sp57_14 202000.000000
Rwpos57_15 in57_15 sp57_15 78000.000000
Rwpos57_16 in57_16 sp57_16 202000.000000
Rwpos57_17 in57_17 sp57_17 78000.000000
Rwpos57_18 in57_18 sp57_18 202000.000000
Rwpos57_19 in57_19 sp57_19 202000.000000
Rwpos57_20 in57_20 sp57_20 202000.000000
Rwpos57_21 in57_21 sp57_21 78000.000000
Rwpos57_22 in57_22 sp57_22 78000.000000
Rwpos57_23 in57_23 sp57_23 78000.000000
Rwpos57_24 in57_24 sp57_24 78000.000000
Rwpos57_25 in57_25 sp57_25 78000.000000
Rwpos57_26 in57_26 sp57_26 202000.000000
Rwpos57_27 in57_27 sp57_27 78000.000000
Rwpos57_28 in57_28 sp57_28 202000.000000
Rwpos57_29 in57_29 sp57_29 202000.000000
Rwpos57_30 in57_30 sp57_30 202000.000000
Rwpos57_31 in57_31 sp57_31 78000.000000
Rwpos57_32 in57_32 sp57_32 78000.000000
Rwpos57_33 in57_33 sp57_33 202000.000000
Rwpos57_34 in57_34 sp57_34 202000.000000
Rwpos57_35 in57_35 sp57_35 202000.000000
Rwpos57_36 in57_36 sp57_36 202000.000000
Rwpos57_37 in57_37 sp57_37 78000.000000
Rwpos57_38 in57_38 sp57_38 202000.000000
Rwpos57_39 in57_39 sp57_39 202000.000000
Rwpos57_40 in57_40 sp57_40 202000.000000
Rwpos57_41 in57_41 sp57_41 202000.000000
Rwpos57_42 in57_42 sp57_42 202000.000000
Rwpos57_43 in57_43 sp57_43 78000.000000
Rwpos57_44 in57_44 sp57_44 78000.000000
Rwpos57_45 in57_45 sp57_45 202000.000000
Rwpos57_46 in57_46 sp57_46 202000.000000
Rwpos57_47 in57_47 sp57_47 202000.000000
Rwpos57_48 in57_48 sp57_48 202000.000000
Rwpos57_49 in57_49 sp57_49 202000.000000
Rwpos57_50 in57_50 sp57_50 202000.000000
Rwpos57_51 in57_51 sp57_51 78000.000000
Rwpos57_52 in57_52 sp57_52 202000.000000
Rwpos57_53 in57_53 sp57_53 78000.000000
Rwpos57_54 in57_54 sp57_54 78000.000000
Rwpos57_55 in57_55 sp57_55 202000.000000
Rwpos57_56 in57_56 sp57_56 78000.000000
Rwpos57_57 in57_57 sp57_57 78000.000000
Rwpos57_58 in57_58 sp57_58 78000.000000
Rwpos57_59 in57_59 sp57_59 202000.000000
Rwpos57_60 in57_60 sp57_60 202000.000000
Rwpos57_61 in57_61 sp57_61 78000.000000
Rwpos57_62 in57_62 sp57_62 78000.000000
Rwpos57_63 in57_63 sp57_63 78000.000000
Rwpos57_64 in57_64 sp57_64 78000.000000
Rwpos57_65 in57_65 sp57_65 78000.000000
Rwpos57_66 in57_66 sp57_66 78000.000000
Rwpos57_67 in57_67 sp57_67 202000.000000
Rwpos57_68 in57_68 sp57_68 78000.000000
Rwpos57_69 in57_69 sp57_69 78000.000000
Rwpos57_70 in57_70 sp57_70 78000.000000
Rwpos57_71 in57_71 sp57_71 202000.000000
Rwpos57_72 in57_72 sp57_72 78000.000000
Rwpos57_73 in57_73 sp57_73 78000.000000
Rwpos57_74 in57_74 sp57_74 78000.000000
Rwpos57_75 in57_75 sp57_75 202000.000000
Rwpos57_76 in57_76 sp57_76 202000.000000
Rwpos57_77 in57_77 sp57_77 202000.000000
Rwpos57_78 in57_78 sp57_78 78000.000000
Rwpos57_79 in57_79 sp57_79 78000.000000
Rwpos57_80 in57_80 sp57_80 78000.000000
Rwpos57_81 in57_81 sp57_81 78000.000000
Rwpos57_82 in57_82 sp57_82 78000.000000
Rwpos57_83 in57_83 sp57_83 202000.000000
Rwpos57_84 in57_84 sp57_84 78000.000000
Rwpos58_1 in58_1 sp58_1 78000.000000
Rwpos58_2 in58_2 sp58_2 78000.000000
Rwpos58_3 in58_3 sp58_3 78000.000000
Rwpos58_4 in58_4 sp58_4 78000.000000
Rwpos58_5 in58_5 sp58_5 202000.000000
Rwpos58_6 in58_6 sp58_6 202000.000000
Rwpos58_7 in58_7 sp58_7 202000.000000
Rwpos58_8 in58_8 sp58_8 202000.000000
Rwpos58_9 in58_9 sp58_9 202000.000000
Rwpos58_10 in58_10 sp58_10 78000.000000
Rwpos58_11 in58_11 sp58_11 202000.000000
Rwpos58_12 in58_12 sp58_12 202000.000000
Rwpos58_13 in58_13 sp58_13 78000.000000
Rwpos58_14 in58_14 sp58_14 78000.000000
Rwpos58_15 in58_15 sp58_15 78000.000000
Rwpos58_16 in58_16 sp58_16 202000.000000
Rwpos58_17 in58_17 sp58_17 78000.000000
Rwpos58_18 in58_18 sp58_18 78000.000000
Rwpos58_19 in58_19 sp58_19 202000.000000
Rwpos58_20 in58_20 sp58_20 78000.000000
Rwpos58_21 in58_21 sp58_21 202000.000000
Rwpos58_22 in58_22 sp58_22 78000.000000
Rwpos58_23 in58_23 sp58_23 78000.000000
Rwpos58_24 in58_24 sp58_24 78000.000000
Rwpos58_25 in58_25 sp58_25 202000.000000
Rwpos58_26 in58_26 sp58_26 202000.000000
Rwpos58_27 in58_27 sp58_27 202000.000000
Rwpos58_28 in58_28 sp58_28 202000.000000
Rwpos58_29 in58_29 sp58_29 78000.000000
Rwpos58_30 in58_30 sp58_30 202000.000000
Rwpos58_31 in58_31 sp58_31 202000.000000
Rwpos58_32 in58_32 sp58_32 78000.000000
Rwpos58_33 in58_33 sp58_33 78000.000000
Rwpos58_34 in58_34 sp58_34 202000.000000
Rwpos58_35 in58_35 sp58_35 78000.000000
Rwpos58_36 in58_36 sp58_36 78000.000000
Rwpos58_37 in58_37 sp58_37 202000.000000
Rwpos58_38 in58_38 sp58_38 202000.000000
Rwpos58_39 in58_39 sp58_39 78000.000000
Rwpos58_40 in58_40 sp58_40 202000.000000
Rwpos58_41 in58_41 sp58_41 202000.000000
Rwpos58_42 in58_42 sp58_42 202000.000000
Rwpos58_43 in58_43 sp58_43 202000.000000
Rwpos58_44 in58_44 sp58_44 202000.000000
Rwpos58_45 in58_45 sp58_45 202000.000000
Rwpos58_46 in58_46 sp58_46 78000.000000
Rwpos58_47 in58_47 sp58_47 78000.000000
Rwpos58_48 in58_48 sp58_48 202000.000000
Rwpos58_49 in58_49 sp58_49 78000.000000
Rwpos58_50 in58_50 sp58_50 78000.000000
Rwpos58_51 in58_51 sp58_51 202000.000000
Rwpos58_52 in58_52 sp58_52 78000.000000
Rwpos58_53 in58_53 sp58_53 78000.000000
Rwpos58_54 in58_54 sp58_54 78000.000000
Rwpos58_55 in58_55 sp58_55 78000.000000
Rwpos58_56 in58_56 sp58_56 202000.000000
Rwpos58_57 in58_57 sp58_57 78000.000000
Rwpos58_58 in58_58 sp58_58 202000.000000
Rwpos58_59 in58_59 sp58_59 202000.000000
Rwpos58_60 in58_60 sp58_60 78000.000000
Rwpos58_61 in58_61 sp58_61 202000.000000
Rwpos58_62 in58_62 sp58_62 78000.000000
Rwpos58_63 in58_63 sp58_63 202000.000000
Rwpos58_64 in58_64 sp58_64 78000.000000
Rwpos58_65 in58_65 sp58_65 202000.000000
Rwpos58_66 in58_66 sp58_66 202000.000000
Rwpos58_67 in58_67 sp58_67 78000.000000
Rwpos58_68 in58_68 sp58_68 202000.000000
Rwpos58_69 in58_69 sp58_69 202000.000000
Rwpos58_70 in58_70 sp58_70 202000.000000
Rwpos58_71 in58_71 sp58_71 202000.000000
Rwpos58_72 in58_72 sp58_72 202000.000000
Rwpos58_73 in58_73 sp58_73 202000.000000
Rwpos58_74 in58_74 sp58_74 78000.000000
Rwpos58_75 in58_75 sp58_75 78000.000000
Rwpos58_76 in58_76 sp58_76 202000.000000
Rwpos58_77 in58_77 sp58_77 202000.000000
Rwpos58_78 in58_78 sp58_78 78000.000000
Rwpos58_79 in58_79 sp58_79 78000.000000
Rwpos58_80 in58_80 sp58_80 202000.000000
Rwpos58_81 in58_81 sp58_81 78000.000000
Rwpos58_82 in58_82 sp58_82 202000.000000
Rwpos58_83 in58_83 sp58_83 78000.000000
Rwpos58_84 in58_84 sp58_84 78000.000000
Rwpos59_1 in59_1 sp59_1 78000.000000
Rwpos59_2 in59_2 sp59_2 202000.000000
Rwpos59_3 in59_3 sp59_3 202000.000000
Rwpos59_4 in59_4 sp59_4 202000.000000
Rwpos59_5 in59_5 sp59_5 202000.000000
Rwpos59_6 in59_6 sp59_6 78000.000000
Rwpos59_7 in59_7 sp59_7 78000.000000
Rwpos59_8 in59_8 sp59_8 202000.000000
Rwpos59_9 in59_9 sp59_9 202000.000000
Rwpos59_10 in59_10 sp59_10 78000.000000
Rwpos59_11 in59_11 sp59_11 78000.000000
Rwpos59_12 in59_12 sp59_12 78000.000000
Rwpos59_13 in59_13 sp59_13 202000.000000
Rwpos59_14 in59_14 sp59_14 202000.000000
Rwpos59_15 in59_15 sp59_15 202000.000000
Rwpos59_16 in59_16 sp59_16 78000.000000
Rwpos59_17 in59_17 sp59_17 78000.000000
Rwpos59_18 in59_18 sp59_18 78000.000000
Rwpos59_19 in59_19 sp59_19 202000.000000
Rwpos59_20 in59_20 sp59_20 202000.000000
Rwpos59_21 in59_21 sp59_21 78000.000000
Rwpos59_22 in59_22 sp59_22 78000.000000
Rwpos59_23 in59_23 sp59_23 78000.000000
Rwpos59_24 in59_24 sp59_24 78000.000000
Rwpos59_25 in59_25 sp59_25 78000.000000
Rwpos59_26 in59_26 sp59_26 202000.000000
Rwpos59_27 in59_27 sp59_27 202000.000000
Rwpos59_28 in59_28 sp59_28 78000.000000
Rwpos59_29 in59_29 sp59_29 78000.000000
Rwpos59_30 in59_30 sp59_30 78000.000000
Rwpos59_31 in59_31 sp59_31 202000.000000
Rwpos59_32 in59_32 sp59_32 78000.000000
Rwpos59_33 in59_33 sp59_33 202000.000000
Rwpos59_34 in59_34 sp59_34 78000.000000
Rwpos59_35 in59_35 sp59_35 78000.000000
Rwpos59_36 in59_36 sp59_36 78000.000000
Rwpos59_37 in59_37 sp59_37 78000.000000
Rwpos59_38 in59_38 sp59_38 202000.000000
Rwpos59_39 in59_39 sp59_39 78000.000000
Rwpos59_40 in59_40 sp59_40 78000.000000
Rwpos59_41 in59_41 sp59_41 78000.000000
Rwpos59_42 in59_42 sp59_42 202000.000000
Rwpos59_43 in59_43 sp59_43 202000.000000
Rwpos59_44 in59_44 sp59_44 202000.000000
Rwpos59_45 in59_45 sp59_45 202000.000000
Rwpos59_46 in59_46 sp59_46 78000.000000
Rwpos59_47 in59_47 sp59_47 78000.000000
Rwpos59_48 in59_48 sp59_48 78000.000000
Rwpos59_49 in59_49 sp59_49 202000.000000
Rwpos59_50 in59_50 sp59_50 202000.000000
Rwpos59_51 in59_51 sp59_51 78000.000000
Rwpos59_52 in59_52 sp59_52 202000.000000
Rwpos59_53 in59_53 sp59_53 78000.000000
Rwpos59_54 in59_54 sp59_54 202000.000000
Rwpos59_55 in59_55 sp59_55 202000.000000
Rwpos59_56 in59_56 sp59_56 202000.000000
Rwpos59_57 in59_57 sp59_57 202000.000000
Rwpos59_58 in59_58 sp59_58 78000.000000
Rwpos59_59 in59_59 sp59_59 78000.000000
Rwpos59_60 in59_60 sp59_60 202000.000000
Rwpos59_61 in59_61 sp59_61 202000.000000
Rwpos59_62 in59_62 sp59_62 78000.000000
Rwpos59_63 in59_63 sp59_63 202000.000000
Rwpos59_64 in59_64 sp59_64 78000.000000
Rwpos59_65 in59_65 sp59_65 78000.000000
Rwpos59_66 in59_66 sp59_66 202000.000000
Rwpos59_67 in59_67 sp59_67 78000.000000
Rwpos59_68 in59_68 sp59_68 78000.000000
Rwpos59_69 in59_69 sp59_69 202000.000000
Rwpos59_70 in59_70 sp59_70 78000.000000
Rwpos59_71 in59_71 sp59_71 202000.000000
Rwpos59_72 in59_72 sp59_72 78000.000000
Rwpos59_73 in59_73 sp59_73 78000.000000
Rwpos59_74 in59_74 sp59_74 78000.000000
Rwpos59_75 in59_75 sp59_75 78000.000000
Rwpos59_76 in59_76 sp59_76 202000.000000
Rwpos59_77 in59_77 sp59_77 78000.000000
Rwpos59_78 in59_78 sp59_78 202000.000000
Rwpos59_79 in59_79 sp59_79 78000.000000
Rwpos59_80 in59_80 sp59_80 78000.000000
Rwpos59_81 in59_81 sp59_81 78000.000000
Rwpos59_82 in59_82 sp59_82 78000.000000
Rwpos59_83 in59_83 sp59_83 202000.000000
Rwpos59_84 in59_84 sp59_84 78000.000000
Rwpos60_1 in60_1 sp60_1 78000.000000
Rwpos60_2 in60_2 sp60_2 78000.000000
Rwpos60_3 in60_3 sp60_3 78000.000000
Rwpos60_4 in60_4 sp60_4 78000.000000
Rwpos60_5 in60_5 sp60_5 202000.000000
Rwpos60_6 in60_6 sp60_6 202000.000000
Rwpos60_7 in60_7 sp60_7 78000.000000
Rwpos60_8 in60_8 sp60_8 78000.000000
Rwpos60_9 in60_9 sp60_9 202000.000000
Rwpos60_10 in60_10 sp60_10 78000.000000
Rwpos60_11 in60_11 sp60_11 78000.000000
Rwpos60_12 in60_12 sp60_12 202000.000000
Rwpos60_13 in60_13 sp60_13 202000.000000
Rwpos60_14 in60_14 sp60_14 202000.000000
Rwpos60_15 in60_15 sp60_15 202000.000000
Rwpos60_16 in60_16 sp60_16 78000.000000
Rwpos60_17 in60_17 sp60_17 202000.000000
Rwpos60_18 in60_18 sp60_18 202000.000000
Rwpos60_19 in60_19 sp60_19 202000.000000
Rwpos60_20 in60_20 sp60_20 78000.000000
Rwpos60_21 in60_21 sp60_21 78000.000000
Rwpos60_22 in60_22 sp60_22 202000.000000
Rwpos60_23 in60_23 sp60_23 78000.000000
Rwpos60_24 in60_24 sp60_24 78000.000000
Rwpos60_25 in60_25 sp60_25 202000.000000
Rwpos60_26 in60_26 sp60_26 78000.000000
Rwpos60_27 in60_27 sp60_27 78000.000000
Rwpos60_28 in60_28 sp60_28 78000.000000
Rwpos60_29 in60_29 sp60_29 78000.000000
Rwpos60_30 in60_30 sp60_30 202000.000000
Rwpos60_31 in60_31 sp60_31 202000.000000
Rwpos60_32 in60_32 sp60_32 202000.000000
Rwpos60_33 in60_33 sp60_33 78000.000000
Rwpos60_34 in60_34 sp60_34 202000.000000
Rwpos60_35 in60_35 sp60_35 78000.000000
Rwpos60_36 in60_36 sp60_36 202000.000000
Rwpos60_37 in60_37 sp60_37 78000.000000
Rwpos60_38 in60_38 sp60_38 202000.000000
Rwpos60_39 in60_39 sp60_39 202000.000000
Rwpos60_40 in60_40 sp60_40 202000.000000
Rwpos60_41 in60_41 sp60_41 202000.000000
Rwpos60_42 in60_42 sp60_42 78000.000000
Rwpos60_43 in60_43 sp60_43 202000.000000
Rwpos60_44 in60_44 sp60_44 78000.000000
Rwpos60_45 in60_45 sp60_45 202000.000000
Rwpos60_46 in60_46 sp60_46 78000.000000
Rwpos60_47 in60_47 sp60_47 202000.000000
Rwpos60_48 in60_48 sp60_48 78000.000000
Rwpos60_49 in60_49 sp60_49 78000.000000
Rwpos60_50 in60_50 sp60_50 202000.000000
Rwpos60_51 in60_51 sp60_51 78000.000000
Rwpos60_52 in60_52 sp60_52 78000.000000
Rwpos60_53 in60_53 sp60_53 202000.000000
Rwpos60_54 in60_54 sp60_54 78000.000000
Rwpos60_55 in60_55 sp60_55 78000.000000
Rwpos60_56 in60_56 sp60_56 202000.000000
Rwpos60_57 in60_57 sp60_57 78000.000000
Rwpos60_58 in60_58 sp60_58 78000.000000
Rwpos60_59 in60_59 sp60_59 202000.000000
Rwpos60_60 in60_60 sp60_60 78000.000000
Rwpos60_61 in60_61 sp60_61 202000.000000
Rwpos60_62 in60_62 sp60_62 78000.000000
Rwpos60_63 in60_63 sp60_63 202000.000000
Rwpos60_64 in60_64 sp60_64 202000.000000
Rwpos60_65 in60_65 sp60_65 78000.000000
Rwpos60_66 in60_66 sp60_66 78000.000000
Rwpos60_67 in60_67 sp60_67 202000.000000
Rwpos60_68 in60_68 sp60_68 202000.000000
Rwpos60_69 in60_69 sp60_69 78000.000000
Rwpos60_70 in60_70 sp60_70 78000.000000
Rwpos60_71 in60_71 sp60_71 202000.000000
Rwpos60_72 in60_72 sp60_72 202000.000000
Rwpos60_73 in60_73 sp60_73 202000.000000
Rwpos60_74 in60_74 sp60_74 202000.000000
Rwpos60_75 in60_75 sp60_75 202000.000000
Rwpos60_76 in60_76 sp60_76 78000.000000
Rwpos60_77 in60_77 sp60_77 202000.000000
Rwpos60_78 in60_78 sp60_78 202000.000000
Rwpos60_79 in60_79 sp60_79 202000.000000
Rwpos60_80 in60_80 sp60_80 202000.000000
Rwpos60_81 in60_81 sp60_81 78000.000000
Rwpos60_82 in60_82 sp60_82 78000.000000
Rwpos60_83 in60_83 sp60_83 202000.000000
Rwpos60_84 in60_84 sp60_84 78000.000000
Rwpos61_1 in61_1 sp61_1 78000.000000
Rwpos61_2 in61_2 sp61_2 202000.000000
Rwpos61_3 in61_3 sp61_3 78000.000000
Rwpos61_4 in61_4 sp61_4 78000.000000
Rwpos61_5 in61_5 sp61_5 78000.000000
Rwpos61_6 in61_6 sp61_6 78000.000000
Rwpos61_7 in61_7 sp61_7 78000.000000
Rwpos61_8 in61_8 sp61_8 202000.000000
Rwpos61_9 in61_9 sp61_9 78000.000000
Rwpos61_10 in61_10 sp61_10 78000.000000
Rwpos61_11 in61_11 sp61_11 202000.000000
Rwpos61_12 in61_12 sp61_12 78000.000000
Rwpos61_13 in61_13 sp61_13 78000.000000
Rwpos61_14 in61_14 sp61_14 78000.000000
Rwpos61_15 in61_15 sp61_15 78000.000000
Rwpos61_16 in61_16 sp61_16 202000.000000
Rwpos61_17 in61_17 sp61_17 78000.000000
Rwpos61_18 in61_18 sp61_18 78000.000000
Rwpos61_19 in61_19 sp61_19 202000.000000
Rwpos61_20 in61_20 sp61_20 202000.000000
Rwpos61_21 in61_21 sp61_21 78000.000000
Rwpos61_22 in61_22 sp61_22 78000.000000
Rwpos61_23 in61_23 sp61_23 202000.000000
Rwpos61_24 in61_24 sp61_24 78000.000000
Rwpos61_25 in61_25 sp61_25 78000.000000
Rwpos61_26 in61_26 sp61_26 202000.000000
Rwpos61_27 in61_27 sp61_27 78000.000000
Rwpos61_28 in61_28 sp61_28 202000.000000
Rwpos61_29 in61_29 sp61_29 78000.000000
Rwpos61_30 in61_30 sp61_30 78000.000000
Rwpos61_31 in61_31 sp61_31 78000.000000
Rwpos61_32 in61_32 sp61_32 202000.000000
Rwpos61_33 in61_33 sp61_33 202000.000000
Rwpos61_34 in61_34 sp61_34 202000.000000
Rwpos61_35 in61_35 sp61_35 202000.000000
Rwpos61_36 in61_36 sp61_36 78000.000000
Rwpos61_37 in61_37 sp61_37 202000.000000
Rwpos61_38 in61_38 sp61_38 202000.000000
Rwpos61_39 in61_39 sp61_39 202000.000000
Rwpos61_40 in61_40 sp61_40 202000.000000
Rwpos61_41 in61_41 sp61_41 78000.000000
Rwpos61_42 in61_42 sp61_42 202000.000000
Rwpos61_43 in61_43 sp61_43 78000.000000
Rwpos61_44 in61_44 sp61_44 78000.000000
Rwpos61_45 in61_45 sp61_45 202000.000000
Rwpos61_46 in61_46 sp61_46 202000.000000
Rwpos61_47 in61_47 sp61_47 78000.000000
Rwpos61_48 in61_48 sp61_48 202000.000000
Rwpos61_49 in61_49 sp61_49 202000.000000
Rwpos61_50 in61_50 sp61_50 78000.000000
Rwpos61_51 in61_51 sp61_51 202000.000000
Rwpos61_52 in61_52 sp61_52 78000.000000
Rwpos61_53 in61_53 sp61_53 202000.000000
Rwpos61_54 in61_54 sp61_54 202000.000000
Rwpos61_55 in61_55 sp61_55 202000.000000
Rwpos61_56 in61_56 sp61_56 78000.000000
Rwpos61_57 in61_57 sp61_57 78000.000000
Rwpos61_58 in61_58 sp61_58 78000.000000
Rwpos61_59 in61_59 sp61_59 78000.000000
Rwpos61_60 in61_60 sp61_60 78000.000000
Rwpos61_61 in61_61 sp61_61 78000.000000
Rwpos61_62 in61_62 sp61_62 78000.000000
Rwpos61_63 in61_63 sp61_63 78000.000000
Rwpos61_64 in61_64 sp61_64 78000.000000
Rwpos61_65 in61_65 sp61_65 202000.000000
Rwpos61_66 in61_66 sp61_66 202000.000000
Rwpos61_67 in61_67 sp61_67 78000.000000
Rwpos61_68 in61_68 sp61_68 78000.000000
Rwpos61_69 in61_69 sp61_69 78000.000000
Rwpos61_70 in61_70 sp61_70 202000.000000
Rwpos61_71 in61_71 sp61_71 78000.000000
Rwpos61_72 in61_72 sp61_72 78000.000000
Rwpos61_73 in61_73 sp61_73 202000.000000
Rwpos61_74 in61_74 sp61_74 78000.000000
Rwpos61_75 in61_75 sp61_75 202000.000000
Rwpos61_76 in61_76 sp61_76 78000.000000
Rwpos61_77 in61_77 sp61_77 202000.000000
Rwpos61_78 in61_78 sp61_78 78000.000000
Rwpos61_79 in61_79 sp61_79 202000.000000
Rwpos61_80 in61_80 sp61_80 202000.000000
Rwpos61_81 in61_81 sp61_81 78000.000000
Rwpos61_82 in61_82 sp61_82 78000.000000
Rwpos61_83 in61_83 sp61_83 78000.000000
Rwpos61_84 in61_84 sp61_84 202000.000000
Rwpos62_1 in62_1 sp62_1 78000.000000
Rwpos62_2 in62_2 sp62_2 202000.000000
Rwpos62_3 in62_3 sp62_3 202000.000000
Rwpos62_4 in62_4 sp62_4 202000.000000
Rwpos62_5 in62_5 sp62_5 202000.000000
Rwpos62_6 in62_6 sp62_6 78000.000000
Rwpos62_7 in62_7 sp62_7 202000.000000
Rwpos62_8 in62_8 sp62_8 202000.000000
Rwpos62_9 in62_9 sp62_9 202000.000000
Rwpos62_10 in62_10 sp62_10 78000.000000
Rwpos62_11 in62_11 sp62_11 78000.000000
Rwpos62_12 in62_12 sp62_12 78000.000000
Rwpos62_13 in62_13 sp62_13 78000.000000
Rwpos62_14 in62_14 sp62_14 202000.000000
Rwpos62_15 in62_15 sp62_15 202000.000000
Rwpos62_16 in62_16 sp62_16 202000.000000
Rwpos62_17 in62_17 sp62_17 78000.000000
Rwpos62_18 in62_18 sp62_18 78000.000000
Rwpos62_19 in62_19 sp62_19 78000.000000
Rwpos62_20 in62_20 sp62_20 78000.000000
Rwpos62_21 in62_21 sp62_21 202000.000000
Rwpos62_22 in62_22 sp62_22 78000.000000
Rwpos62_23 in62_23 sp62_23 78000.000000
Rwpos62_24 in62_24 sp62_24 202000.000000
Rwpos62_25 in62_25 sp62_25 78000.000000
Rwpos62_26 in62_26 sp62_26 78000.000000
Rwpos62_27 in62_27 sp62_27 78000.000000
Rwpos62_28 in62_28 sp62_28 78000.000000
Rwpos62_29 in62_29 sp62_29 202000.000000
Rwpos62_30 in62_30 sp62_30 78000.000000
Rwpos62_31 in62_31 sp62_31 78000.000000
Rwpos62_32 in62_32 sp62_32 78000.000000
Rwpos62_33 in62_33 sp62_33 78000.000000
Rwpos62_34 in62_34 sp62_34 202000.000000
Rwpos62_35 in62_35 sp62_35 202000.000000
Rwpos62_36 in62_36 sp62_36 202000.000000
Rwpos62_37 in62_37 sp62_37 78000.000000
Rwpos62_38 in62_38 sp62_38 202000.000000
Rwpos62_39 in62_39 sp62_39 202000.000000
Rwpos62_40 in62_40 sp62_40 78000.000000
Rwpos62_41 in62_41 sp62_41 202000.000000
Rwpos62_42 in62_42 sp62_42 202000.000000
Rwpos62_43 in62_43 sp62_43 202000.000000
Rwpos62_44 in62_44 sp62_44 202000.000000
Rwpos62_45 in62_45 sp62_45 78000.000000
Rwpos62_46 in62_46 sp62_46 202000.000000
Rwpos62_47 in62_47 sp62_47 202000.000000
Rwpos62_48 in62_48 sp62_48 78000.000000
Rwpos62_49 in62_49 sp62_49 202000.000000
Rwpos62_50 in62_50 sp62_50 202000.000000
Rwpos62_51 in62_51 sp62_51 78000.000000
Rwpos62_52 in62_52 sp62_52 202000.000000
Rwpos62_53 in62_53 sp62_53 202000.000000
Rwpos62_54 in62_54 sp62_54 78000.000000
Rwpos62_55 in62_55 sp62_55 78000.000000
Rwpos62_56 in62_56 sp62_56 78000.000000
Rwpos62_57 in62_57 sp62_57 202000.000000
Rwpos62_58 in62_58 sp62_58 78000.000000
Rwpos62_59 in62_59 sp62_59 202000.000000
Rwpos62_60 in62_60 sp62_60 202000.000000
Rwpos62_61 in62_61 sp62_61 78000.000000
Rwpos62_62 in62_62 sp62_62 78000.000000
Rwpos62_63 in62_63 sp62_63 78000.000000
Rwpos62_64 in62_64 sp62_64 78000.000000
Rwpos62_65 in62_65 sp62_65 202000.000000
Rwpos62_66 in62_66 sp62_66 78000.000000
Rwpos62_67 in62_67 sp62_67 78000.000000
Rwpos62_68 in62_68 sp62_68 202000.000000
Rwpos62_69 in62_69 sp62_69 78000.000000
Rwpos62_70 in62_70 sp62_70 78000.000000
Rwpos62_71 in62_71 sp62_71 78000.000000
Rwpos62_72 in62_72 sp62_72 202000.000000
Rwpos62_73 in62_73 sp62_73 78000.000000
Rwpos62_74 in62_74 sp62_74 202000.000000
Rwpos62_75 in62_75 sp62_75 78000.000000
Rwpos62_76 in62_76 sp62_76 202000.000000
Rwpos62_77 in62_77 sp62_77 78000.000000
Rwpos62_78 in62_78 sp62_78 202000.000000
Rwpos62_79 in62_79 sp62_79 78000.000000
Rwpos62_80 in62_80 sp62_80 78000.000000
Rwpos62_81 in62_81 sp62_81 78000.000000
Rwpos62_82 in62_82 sp62_82 78000.000000
Rwpos62_83 in62_83 sp62_83 78000.000000
Rwpos62_84 in62_84 sp62_84 78000.000000
Rwpos63_1 in63_1 sp63_1 202000.000000
Rwpos63_2 in63_2 sp63_2 202000.000000
Rwpos63_3 in63_3 sp63_3 202000.000000
Rwpos63_4 in63_4 sp63_4 202000.000000
Rwpos63_5 in63_5 sp63_5 202000.000000
Rwpos63_6 in63_6 sp63_6 78000.000000
Rwpos63_7 in63_7 sp63_7 78000.000000
Rwpos63_8 in63_8 sp63_8 202000.000000
Rwpos63_9 in63_9 sp63_9 202000.000000
Rwpos63_10 in63_10 sp63_10 78000.000000
Rwpos63_11 in63_11 sp63_11 202000.000000
Rwpos63_12 in63_12 sp63_12 78000.000000
Rwpos63_13 in63_13 sp63_13 202000.000000
Rwpos63_14 in63_14 sp63_14 78000.000000
Rwpos63_15 in63_15 sp63_15 78000.000000
Rwpos63_16 in63_16 sp63_16 78000.000000
Rwpos63_17 in63_17 sp63_17 202000.000000
Rwpos63_18 in63_18 sp63_18 202000.000000
Rwpos63_19 in63_19 sp63_19 78000.000000
Rwpos63_20 in63_20 sp63_20 78000.000000
Rwpos63_21 in63_21 sp63_21 78000.000000
Rwpos63_22 in63_22 sp63_22 202000.000000
Rwpos63_23 in63_23 sp63_23 202000.000000
Rwpos63_24 in63_24 sp63_24 78000.000000
Rwpos63_25 in63_25 sp63_25 78000.000000
Rwpos63_26 in63_26 sp63_26 78000.000000
Rwpos63_27 in63_27 sp63_27 78000.000000
Rwpos63_28 in63_28 sp63_28 78000.000000
Rwpos63_29 in63_29 sp63_29 78000.000000
Rwpos63_30 in63_30 sp63_30 78000.000000
Rwpos63_31 in63_31 sp63_31 202000.000000
Rwpos63_32 in63_32 sp63_32 78000.000000
Rwpos63_33 in63_33 sp63_33 202000.000000
Rwpos63_34 in63_34 sp63_34 78000.000000
Rwpos63_35 in63_35 sp63_35 202000.000000
Rwpos63_36 in63_36 sp63_36 78000.000000
Rwpos63_37 in63_37 sp63_37 78000.000000
Rwpos63_38 in63_38 sp63_38 78000.000000
Rwpos63_39 in63_39 sp63_39 78000.000000
Rwpos63_40 in63_40 sp63_40 78000.000000
Rwpos63_41 in63_41 sp63_41 202000.000000
Rwpos63_42 in63_42 sp63_42 202000.000000
Rwpos63_43 in63_43 sp63_43 78000.000000
Rwpos63_44 in63_44 sp63_44 78000.000000
Rwpos63_45 in63_45 sp63_45 78000.000000
Rwpos63_46 in63_46 sp63_46 78000.000000
Rwpos63_47 in63_47 sp63_47 78000.000000
Rwpos63_48 in63_48 sp63_48 78000.000000
Rwpos63_49 in63_49 sp63_49 78000.000000
Rwpos63_50 in63_50 sp63_50 78000.000000
Rwpos63_51 in63_51 sp63_51 78000.000000
Rwpos63_52 in63_52 sp63_52 78000.000000
Rwpos63_53 in63_53 sp63_53 202000.000000
Rwpos63_54 in63_54 sp63_54 202000.000000
Rwpos63_55 in63_55 sp63_55 202000.000000
Rwpos63_56 in63_56 sp63_56 202000.000000
Rwpos63_57 in63_57 sp63_57 202000.000000
Rwpos63_58 in63_58 sp63_58 202000.000000
Rwpos63_59 in63_59 sp63_59 202000.000000
Rwpos63_60 in63_60 sp63_60 78000.000000
Rwpos63_61 in63_61 sp63_61 202000.000000
Rwpos63_62 in63_62 sp63_62 202000.000000
Rwpos63_63 in63_63 sp63_63 78000.000000
Rwpos63_64 in63_64 sp63_64 202000.000000
Rwpos63_65 in63_65 sp63_65 202000.000000
Rwpos63_66 in63_66 sp63_66 78000.000000
Rwpos63_67 in63_67 sp63_67 78000.000000
Rwpos63_68 in63_68 sp63_68 78000.000000
Rwpos63_69 in63_69 sp63_69 202000.000000
Rwpos63_70 in63_70 sp63_70 78000.000000
Rwpos63_71 in63_71 sp63_71 202000.000000
Rwpos63_72 in63_72 sp63_72 78000.000000
Rwpos63_73 in63_73 sp63_73 202000.000000
Rwpos63_74 in63_74 sp63_74 202000.000000
Rwpos63_75 in63_75 sp63_75 202000.000000
Rwpos63_76 in63_76 sp63_76 78000.000000
Rwpos63_77 in63_77 sp63_77 202000.000000
Rwpos63_78 in63_78 sp63_78 202000.000000
Rwpos63_79 in63_79 sp63_79 78000.000000
Rwpos63_80 in63_80 sp63_80 202000.000000
Rwpos63_81 in63_81 sp63_81 202000.000000
Rwpos63_82 in63_82 sp63_82 78000.000000
Rwpos63_83 in63_83 sp63_83 202000.000000
Rwpos63_84 in63_84 sp63_84 202000.000000
Rwpos64_1 in64_1 sp64_1 78000.000000
Rwpos64_2 in64_2 sp64_2 78000.000000
Rwpos64_3 in64_3 sp64_3 78000.000000
Rwpos64_4 in64_4 sp64_4 78000.000000
Rwpos64_5 in64_5 sp64_5 202000.000000
Rwpos64_6 in64_6 sp64_6 78000.000000
Rwpos64_7 in64_7 sp64_7 78000.000000
Rwpos64_8 in64_8 sp64_8 78000.000000
Rwpos64_9 in64_9 sp64_9 78000.000000
Rwpos64_10 in64_10 sp64_10 78000.000000
Rwpos64_11 in64_11 sp64_11 202000.000000
Rwpos64_12 in64_12 sp64_12 202000.000000
Rwpos64_13 in64_13 sp64_13 202000.000000
Rwpos64_14 in64_14 sp64_14 78000.000000
Rwpos64_15 in64_15 sp64_15 78000.000000
Rwpos64_16 in64_16 sp64_16 78000.000000
Rwpos64_17 in64_17 sp64_17 78000.000000
Rwpos64_18 in64_18 sp64_18 202000.000000
Rwpos64_19 in64_19 sp64_19 202000.000000
Rwpos64_20 in64_20 sp64_20 202000.000000
Rwpos64_21 in64_21 sp64_21 78000.000000
Rwpos64_22 in64_22 sp64_22 78000.000000
Rwpos64_23 in64_23 sp64_23 202000.000000
Rwpos64_24 in64_24 sp64_24 202000.000000
Rwpos64_25 in64_25 sp64_25 202000.000000
Rwpos64_26 in64_26 sp64_26 78000.000000
Rwpos64_27 in64_27 sp64_27 78000.000000
Rwpos64_28 in64_28 sp64_28 202000.000000
Rwpos64_29 in64_29 sp64_29 202000.000000
Rwpos64_30 in64_30 sp64_30 78000.000000
Rwpos64_31 in64_31 sp64_31 78000.000000
Rwpos64_32 in64_32 sp64_32 78000.000000
Rwpos64_33 in64_33 sp64_33 78000.000000
Rwpos64_34 in64_34 sp64_34 202000.000000
Rwpos64_35 in64_35 sp64_35 78000.000000
Rwpos64_36 in64_36 sp64_36 202000.000000
Rwpos64_37 in64_37 sp64_37 202000.000000
Rwpos64_38 in64_38 sp64_38 78000.000000
Rwpos64_39 in64_39 sp64_39 202000.000000
Rwpos64_40 in64_40 sp64_40 202000.000000
Rwpos64_41 in64_41 sp64_41 78000.000000
Rwpos64_42 in64_42 sp64_42 78000.000000
Rwpos64_43 in64_43 sp64_43 202000.000000
Rwpos64_44 in64_44 sp64_44 78000.000000
Rwpos64_45 in64_45 sp64_45 78000.000000
Rwpos64_46 in64_46 sp64_46 78000.000000
Rwpos64_47 in64_47 sp64_47 78000.000000
Rwpos64_48 in64_48 sp64_48 78000.000000
Rwpos64_49 in64_49 sp64_49 202000.000000
Rwpos64_50 in64_50 sp64_50 78000.000000
Rwpos64_51 in64_51 sp64_51 78000.000000
Rwpos64_52 in64_52 sp64_52 78000.000000
Rwpos64_53 in64_53 sp64_53 202000.000000
Rwpos64_54 in64_54 sp64_54 202000.000000
Rwpos64_55 in64_55 sp64_55 202000.000000
Rwpos64_56 in64_56 sp64_56 202000.000000
Rwpos64_57 in64_57 sp64_57 78000.000000
Rwpos64_58 in64_58 sp64_58 78000.000000
Rwpos64_59 in64_59 sp64_59 202000.000000
Rwpos64_60 in64_60 sp64_60 78000.000000
Rwpos64_61 in64_61 sp64_61 78000.000000
Rwpos64_62 in64_62 sp64_62 202000.000000
Rwpos64_63 in64_63 sp64_63 202000.000000
Rwpos64_64 in64_64 sp64_64 78000.000000
Rwpos64_65 in64_65 sp64_65 202000.000000
Rwpos64_66 in64_66 sp64_66 202000.000000
Rwpos64_67 in64_67 sp64_67 78000.000000
Rwpos64_68 in64_68 sp64_68 202000.000000
Rwpos64_69 in64_69 sp64_69 202000.000000
Rwpos64_70 in64_70 sp64_70 78000.000000
Rwpos64_71 in64_71 sp64_71 202000.000000
Rwpos64_72 in64_72 sp64_72 78000.000000
Rwpos64_73 in64_73 sp64_73 78000.000000
Rwpos64_74 in64_74 sp64_74 78000.000000
Rwpos64_75 in64_75 sp64_75 78000.000000
Rwpos64_76 in64_76 sp64_76 78000.000000
Rwpos64_77 in64_77 sp64_77 202000.000000
Rwpos64_78 in64_78 sp64_78 78000.000000
Rwpos64_79 in64_79 sp64_79 202000.000000
Rwpos64_80 in64_80 sp64_80 202000.000000
Rwpos64_81 in64_81 sp64_81 78000.000000
Rwpos64_82 in64_82 sp64_82 202000.000000
Rwpos64_83 in64_83 sp64_83 78000.000000
Rwpos64_84 in64_84 sp64_84 78000.000000
Rwpos65_1 in65_1 sp65_1 78000.000000
Rwpos65_2 in65_2 sp65_2 202000.000000
Rwpos65_3 in65_3 sp65_3 78000.000000
Rwpos65_4 in65_4 sp65_4 78000.000000
Rwpos65_5 in65_5 sp65_5 78000.000000
Rwpos65_6 in65_6 sp65_6 202000.000000
Rwpos65_7 in65_7 sp65_7 202000.000000
Rwpos65_8 in65_8 sp65_8 78000.000000
Rwpos65_9 in65_9 sp65_9 202000.000000
Rwpos65_10 in65_10 sp65_10 202000.000000
Rwpos65_11 in65_11 sp65_11 202000.000000
Rwpos65_12 in65_12 sp65_12 202000.000000
Rwpos65_13 in65_13 sp65_13 78000.000000
Rwpos65_14 in65_14 sp65_14 78000.000000
Rwpos65_15 in65_15 sp65_15 202000.000000
Rwpos65_16 in65_16 sp65_16 202000.000000
Rwpos65_17 in65_17 sp65_17 202000.000000
Rwpos65_18 in65_18 sp65_18 78000.000000
Rwpos65_19 in65_19 sp65_19 78000.000000
Rwpos65_20 in65_20 sp65_20 78000.000000
Rwpos65_21 in65_21 sp65_21 202000.000000
Rwpos65_22 in65_22 sp65_22 202000.000000
Rwpos65_23 in65_23 sp65_23 78000.000000
Rwpos65_24 in65_24 sp65_24 202000.000000
Rwpos65_25 in65_25 sp65_25 78000.000000
Rwpos65_26 in65_26 sp65_26 78000.000000
Rwpos65_27 in65_27 sp65_27 78000.000000
Rwpos65_28 in65_28 sp65_28 78000.000000
Rwpos65_29 in65_29 sp65_29 202000.000000
Rwpos65_30 in65_30 sp65_30 78000.000000
Rwpos65_31 in65_31 sp65_31 78000.000000
Rwpos65_32 in65_32 sp65_32 78000.000000
Rwpos65_33 in65_33 sp65_33 78000.000000
Rwpos65_34 in65_34 sp65_34 202000.000000
Rwpos65_35 in65_35 sp65_35 78000.000000
Rwpos65_36 in65_36 sp65_36 202000.000000
Rwpos65_37 in65_37 sp65_37 78000.000000
Rwpos65_38 in65_38 sp65_38 78000.000000
Rwpos65_39 in65_39 sp65_39 202000.000000
Rwpos65_40 in65_40 sp65_40 78000.000000
Rwpos65_41 in65_41 sp65_41 202000.000000
Rwpos65_42 in65_42 sp65_42 78000.000000
Rwpos65_43 in65_43 sp65_43 78000.000000
Rwpos65_44 in65_44 sp65_44 202000.000000
Rwpos65_45 in65_45 sp65_45 78000.000000
Rwpos65_46 in65_46 sp65_46 78000.000000
Rwpos65_47 in65_47 sp65_47 202000.000000
Rwpos65_48 in65_48 sp65_48 202000.000000
Rwpos65_49 in65_49 sp65_49 78000.000000
Rwpos65_50 in65_50 sp65_50 78000.000000
Rwpos65_51 in65_51 sp65_51 78000.000000
Rwpos65_52 in65_52 sp65_52 78000.000000
Rwpos65_53 in65_53 sp65_53 78000.000000
Rwpos65_54 in65_54 sp65_54 78000.000000
Rwpos65_55 in65_55 sp65_55 202000.000000
Rwpos65_56 in65_56 sp65_56 78000.000000
Rwpos65_57 in65_57 sp65_57 202000.000000
Rwpos65_58 in65_58 sp65_58 202000.000000
Rwpos65_59 in65_59 sp65_59 78000.000000
Rwpos65_60 in65_60 sp65_60 202000.000000
Rwpos65_61 in65_61 sp65_61 202000.000000
Rwpos65_62 in65_62 sp65_62 78000.000000
Rwpos65_63 in65_63 sp65_63 202000.000000
Rwpos65_64 in65_64 sp65_64 202000.000000
Rwpos65_65 in65_65 sp65_65 202000.000000
Rwpos65_66 in65_66 sp65_66 78000.000000
Rwpos65_67 in65_67 sp65_67 78000.000000
Rwpos65_68 in65_68 sp65_68 202000.000000
Rwpos65_69 in65_69 sp65_69 202000.000000
Rwpos65_70 in65_70 sp65_70 202000.000000
Rwpos65_71 in65_71 sp65_71 202000.000000
Rwpos65_72 in65_72 sp65_72 202000.000000
Rwpos65_73 in65_73 sp65_73 202000.000000
Rwpos65_74 in65_74 sp65_74 78000.000000
Rwpos65_75 in65_75 sp65_75 78000.000000
Rwpos65_76 in65_76 sp65_76 202000.000000
Rwpos65_77 in65_77 sp65_77 78000.000000
Rwpos65_78 in65_78 sp65_78 78000.000000
Rwpos65_79 in65_79 sp65_79 202000.000000
Rwpos65_80 in65_80 sp65_80 78000.000000
Rwpos65_81 in65_81 sp65_81 202000.000000
Rwpos65_82 in65_82 sp65_82 202000.000000
Rwpos65_83 in65_83 sp65_83 78000.000000
Rwpos65_84 in65_84 sp65_84 78000.000000
Rwpos66_1 in66_1 sp66_1 78000.000000
Rwpos66_2 in66_2 sp66_2 202000.000000
Rwpos66_3 in66_3 sp66_3 78000.000000
Rwpos66_4 in66_4 sp66_4 202000.000000
Rwpos66_5 in66_5 sp66_5 78000.000000
Rwpos66_6 in66_6 sp66_6 202000.000000
Rwpos66_7 in66_7 sp66_7 78000.000000
Rwpos66_8 in66_8 sp66_8 202000.000000
Rwpos66_9 in66_9 sp66_9 78000.000000
Rwpos66_10 in66_10 sp66_10 202000.000000
Rwpos66_11 in66_11 sp66_11 202000.000000
Rwpos66_12 in66_12 sp66_12 202000.000000
Rwpos66_13 in66_13 sp66_13 202000.000000
Rwpos66_14 in66_14 sp66_14 78000.000000
Rwpos66_15 in66_15 sp66_15 78000.000000
Rwpos66_16 in66_16 sp66_16 78000.000000
Rwpos66_17 in66_17 sp66_17 202000.000000
Rwpos66_18 in66_18 sp66_18 202000.000000
Rwpos66_19 in66_19 sp66_19 202000.000000
Rwpos66_20 in66_20 sp66_20 78000.000000
Rwpos66_21 in66_21 sp66_21 78000.000000
Rwpos66_22 in66_22 sp66_22 202000.000000
Rwpos66_23 in66_23 sp66_23 202000.000000
Rwpos66_24 in66_24 sp66_24 78000.000000
Rwpos66_25 in66_25 sp66_25 202000.000000
Rwpos66_26 in66_26 sp66_26 78000.000000
Rwpos66_27 in66_27 sp66_27 202000.000000
Rwpos66_28 in66_28 sp66_28 78000.000000
Rwpos66_29 in66_29 sp66_29 78000.000000
Rwpos66_30 in66_30 sp66_30 78000.000000
Rwpos66_31 in66_31 sp66_31 202000.000000
Rwpos66_32 in66_32 sp66_32 202000.000000
Rwpos66_33 in66_33 sp66_33 78000.000000
Rwpos66_34 in66_34 sp66_34 202000.000000
Rwpos66_35 in66_35 sp66_35 78000.000000
Rwpos66_36 in66_36 sp66_36 202000.000000
Rwpos66_37 in66_37 sp66_37 78000.000000
Rwpos66_38 in66_38 sp66_38 202000.000000
Rwpos66_39 in66_39 sp66_39 202000.000000
Rwpos66_40 in66_40 sp66_40 202000.000000
Rwpos66_41 in66_41 sp66_41 78000.000000
Rwpos66_42 in66_42 sp66_42 78000.000000
Rwpos66_43 in66_43 sp66_43 78000.000000
Rwpos66_44 in66_44 sp66_44 78000.000000
Rwpos66_45 in66_45 sp66_45 202000.000000
Rwpos66_46 in66_46 sp66_46 202000.000000
Rwpos66_47 in66_47 sp66_47 202000.000000
Rwpos66_48 in66_48 sp66_48 202000.000000
Rwpos66_49 in66_49 sp66_49 78000.000000
Rwpos66_50 in66_50 sp66_50 78000.000000
Rwpos66_51 in66_51 sp66_51 78000.000000
Rwpos66_52 in66_52 sp66_52 78000.000000
Rwpos66_53 in66_53 sp66_53 202000.000000
Rwpos66_54 in66_54 sp66_54 78000.000000
Rwpos66_55 in66_55 sp66_55 78000.000000
Rwpos66_56 in66_56 sp66_56 202000.000000
Rwpos66_57 in66_57 sp66_57 78000.000000
Rwpos66_58 in66_58 sp66_58 202000.000000
Rwpos66_59 in66_59 sp66_59 78000.000000
Rwpos66_60 in66_60 sp66_60 202000.000000
Rwpos66_61 in66_61 sp66_61 78000.000000
Rwpos66_62 in66_62 sp66_62 78000.000000
Rwpos66_63 in66_63 sp66_63 78000.000000
Rwpos66_64 in66_64 sp66_64 202000.000000
Rwpos66_65 in66_65 sp66_65 78000.000000
Rwpos66_66 in66_66 sp66_66 78000.000000
Rwpos66_67 in66_67 sp66_67 202000.000000
Rwpos66_68 in66_68 sp66_68 202000.000000
Rwpos66_69 in66_69 sp66_69 202000.000000
Rwpos66_70 in66_70 sp66_70 78000.000000
Rwpos66_71 in66_71 sp66_71 202000.000000
Rwpos66_72 in66_72 sp66_72 78000.000000
Rwpos66_73 in66_73 sp66_73 202000.000000
Rwpos66_74 in66_74 sp66_74 202000.000000
Rwpos66_75 in66_75 sp66_75 202000.000000
Rwpos66_76 in66_76 sp66_76 78000.000000
Rwpos66_77 in66_77 sp66_77 202000.000000
Rwpos66_78 in66_78 sp66_78 202000.000000
Rwpos66_79 in66_79 sp66_79 202000.000000
Rwpos66_80 in66_80 sp66_80 78000.000000
Rwpos66_81 in66_81 sp66_81 78000.000000
Rwpos66_82 in66_82 sp66_82 78000.000000
Rwpos66_83 in66_83 sp66_83 202000.000000
Rwpos66_84 in66_84 sp66_84 78000.000000
Rwpos67_1 in67_1 sp67_1 202000.000000
Rwpos67_2 in67_2 sp67_2 202000.000000
Rwpos67_3 in67_3 sp67_3 78000.000000
Rwpos67_4 in67_4 sp67_4 202000.000000
Rwpos67_5 in67_5 sp67_5 78000.000000
Rwpos67_6 in67_6 sp67_6 202000.000000
Rwpos67_7 in67_7 sp67_7 78000.000000
Rwpos67_8 in67_8 sp67_8 202000.000000
Rwpos67_9 in67_9 sp67_9 202000.000000
Rwpos67_10 in67_10 sp67_10 78000.000000
Rwpos67_11 in67_11 sp67_11 202000.000000
Rwpos67_12 in67_12 sp67_12 202000.000000
Rwpos67_13 in67_13 sp67_13 202000.000000
Rwpos67_14 in67_14 sp67_14 202000.000000
Rwpos67_15 in67_15 sp67_15 202000.000000
Rwpos67_16 in67_16 sp67_16 78000.000000
Rwpos67_17 in67_17 sp67_17 78000.000000
Rwpos67_18 in67_18 sp67_18 202000.000000
Rwpos67_19 in67_19 sp67_19 78000.000000
Rwpos67_20 in67_20 sp67_20 202000.000000
Rwpos67_21 in67_21 sp67_21 78000.000000
Rwpos67_22 in67_22 sp67_22 78000.000000
Rwpos67_23 in67_23 sp67_23 78000.000000
Rwpos67_24 in67_24 sp67_24 78000.000000
Rwpos67_25 in67_25 sp67_25 202000.000000
Rwpos67_26 in67_26 sp67_26 202000.000000
Rwpos67_27 in67_27 sp67_27 78000.000000
Rwpos67_28 in67_28 sp67_28 78000.000000
Rwpos67_29 in67_29 sp67_29 78000.000000
Rwpos67_30 in67_30 sp67_30 78000.000000
Rwpos67_31 in67_31 sp67_31 78000.000000
Rwpos67_32 in67_32 sp67_32 78000.000000
Rwpos67_33 in67_33 sp67_33 78000.000000
Rwpos67_34 in67_34 sp67_34 202000.000000
Rwpos67_35 in67_35 sp67_35 202000.000000
Rwpos67_36 in67_36 sp67_36 202000.000000
Rwpos67_37 in67_37 sp67_37 78000.000000
Rwpos67_38 in67_38 sp67_38 78000.000000
Rwpos67_39 in67_39 sp67_39 202000.000000
Rwpos67_40 in67_40 sp67_40 202000.000000
Rwpos67_41 in67_41 sp67_41 202000.000000
Rwpos67_42 in67_42 sp67_42 202000.000000
Rwpos67_43 in67_43 sp67_43 202000.000000
Rwpos67_44 in67_44 sp67_44 78000.000000
Rwpos67_45 in67_45 sp67_45 78000.000000
Rwpos67_46 in67_46 sp67_46 78000.000000
Rwpos67_47 in67_47 sp67_47 202000.000000
Rwpos67_48 in67_48 sp67_48 78000.000000
Rwpos67_49 in67_49 sp67_49 202000.000000
Rwpos67_50 in67_50 sp67_50 202000.000000
Rwpos67_51 in67_51 sp67_51 78000.000000
Rwpos67_52 in67_52 sp67_52 202000.000000
Rwpos67_53 in67_53 sp67_53 202000.000000
Rwpos67_54 in67_54 sp67_54 78000.000000
Rwpos67_55 in67_55 sp67_55 78000.000000
Rwpos67_56 in67_56 sp67_56 202000.000000
Rwpos67_57 in67_57 sp67_57 78000.000000
Rwpos67_58 in67_58 sp67_58 78000.000000
Rwpos67_59 in67_59 sp67_59 78000.000000
Rwpos67_60 in67_60 sp67_60 202000.000000
Rwpos67_61 in67_61 sp67_61 78000.000000
Rwpos67_62 in67_62 sp67_62 78000.000000
Rwpos67_63 in67_63 sp67_63 202000.000000
Rwpos67_64 in67_64 sp67_64 78000.000000
Rwpos67_65 in67_65 sp67_65 202000.000000
Rwpos67_66 in67_66 sp67_66 202000.000000
Rwpos67_67 in67_67 sp67_67 78000.000000
Rwpos67_68 in67_68 sp67_68 202000.000000
Rwpos67_69 in67_69 sp67_69 202000.000000
Rwpos67_70 in67_70 sp67_70 78000.000000
Rwpos67_71 in67_71 sp67_71 202000.000000
Rwpos67_72 in67_72 sp67_72 78000.000000
Rwpos67_73 in67_73 sp67_73 78000.000000
Rwpos67_74 in67_74 sp67_74 78000.000000
Rwpos67_75 in67_75 sp67_75 78000.000000
Rwpos67_76 in67_76 sp67_76 202000.000000
Rwpos67_77 in67_77 sp67_77 78000.000000
Rwpos67_78 in67_78 sp67_78 78000.000000
Rwpos67_79 in67_79 sp67_79 202000.000000
Rwpos67_80 in67_80 sp67_80 78000.000000
Rwpos67_81 in67_81 sp67_81 78000.000000
Rwpos67_82 in67_82 sp67_82 202000.000000
Rwpos67_83 in67_83 sp67_83 78000.000000
Rwpos67_84 in67_84 sp67_84 202000.000000
Rwpos68_1 in68_1 sp68_1 78000.000000
Rwpos68_2 in68_2 sp68_2 78000.000000
Rwpos68_3 in68_3 sp68_3 78000.000000
Rwpos68_4 in68_4 sp68_4 202000.000000
Rwpos68_5 in68_5 sp68_5 202000.000000
Rwpos68_6 in68_6 sp68_6 78000.000000
Rwpos68_7 in68_7 sp68_7 202000.000000
Rwpos68_8 in68_8 sp68_8 202000.000000
Rwpos68_9 in68_9 sp68_9 202000.000000
Rwpos68_10 in68_10 sp68_10 78000.000000
Rwpos68_11 in68_11 sp68_11 202000.000000
Rwpos68_12 in68_12 sp68_12 202000.000000
Rwpos68_13 in68_13 sp68_13 202000.000000
Rwpos68_14 in68_14 sp68_14 78000.000000
Rwpos68_15 in68_15 sp68_15 202000.000000
Rwpos68_16 in68_16 sp68_16 202000.000000
Rwpos68_17 in68_17 sp68_17 202000.000000
Rwpos68_18 in68_18 sp68_18 78000.000000
Rwpos68_19 in68_19 sp68_19 78000.000000
Rwpos68_20 in68_20 sp68_20 78000.000000
Rwpos68_21 in68_21 sp68_21 78000.000000
Rwpos68_22 in68_22 sp68_22 78000.000000
Rwpos68_23 in68_23 sp68_23 202000.000000
Rwpos68_24 in68_24 sp68_24 78000.000000
Rwpos68_25 in68_25 sp68_25 202000.000000
Rwpos68_26 in68_26 sp68_26 78000.000000
Rwpos68_27 in68_27 sp68_27 78000.000000
Rwpos68_28 in68_28 sp68_28 78000.000000
Rwpos68_29 in68_29 sp68_29 202000.000000
Rwpos68_30 in68_30 sp68_30 202000.000000
Rwpos68_31 in68_31 sp68_31 202000.000000
Rwpos68_32 in68_32 sp68_32 78000.000000
Rwpos68_33 in68_33 sp68_33 78000.000000
Rwpos68_34 in68_34 sp68_34 202000.000000
Rwpos68_35 in68_35 sp68_35 78000.000000
Rwpos68_36 in68_36 sp68_36 78000.000000
Rwpos68_37 in68_37 sp68_37 78000.000000
Rwpos68_38 in68_38 sp68_38 78000.000000
Rwpos68_39 in68_39 sp68_39 202000.000000
Rwpos68_40 in68_40 sp68_40 202000.000000
Rwpos68_41 in68_41 sp68_41 202000.000000
Rwpos68_42 in68_42 sp68_42 78000.000000
Rwpos68_43 in68_43 sp68_43 78000.000000
Rwpos68_44 in68_44 sp68_44 78000.000000
Rwpos68_45 in68_45 sp68_45 78000.000000
Rwpos68_46 in68_46 sp68_46 202000.000000
Rwpos68_47 in68_47 sp68_47 202000.000000
Rwpos68_48 in68_48 sp68_48 202000.000000
Rwpos68_49 in68_49 sp68_49 202000.000000
Rwpos68_50 in68_50 sp68_50 78000.000000
Rwpos68_51 in68_51 sp68_51 78000.000000
Rwpos68_52 in68_52 sp68_52 78000.000000
Rwpos68_53 in68_53 sp68_53 202000.000000
Rwpos68_54 in68_54 sp68_54 202000.000000
Rwpos68_55 in68_55 sp68_55 202000.000000
Rwpos68_56 in68_56 sp68_56 202000.000000
Rwpos68_57 in68_57 sp68_57 78000.000000
Rwpos68_58 in68_58 sp68_58 202000.000000
Rwpos68_59 in68_59 sp68_59 78000.000000
Rwpos68_60 in68_60 sp68_60 202000.000000
Rwpos68_61 in68_61 sp68_61 78000.000000
Rwpos68_62 in68_62 sp68_62 202000.000000
Rwpos68_63 in68_63 sp68_63 202000.000000
Rwpos68_64 in68_64 sp68_64 78000.000000
Rwpos68_65 in68_65 sp68_65 202000.000000
Rwpos68_66 in68_66 sp68_66 202000.000000
Rwpos68_67 in68_67 sp68_67 78000.000000
Rwpos68_68 in68_68 sp68_68 202000.000000
Rwpos68_69 in68_69 sp68_69 202000.000000
Rwpos68_70 in68_70 sp68_70 202000.000000
Rwpos68_71 in68_71 sp68_71 202000.000000
Rwpos68_72 in68_72 sp68_72 78000.000000
Rwpos68_73 in68_73 sp68_73 202000.000000
Rwpos68_74 in68_74 sp68_74 202000.000000
Rwpos68_75 in68_75 sp68_75 78000.000000
Rwpos68_76 in68_76 sp68_76 202000.000000
Rwpos68_77 in68_77 sp68_77 78000.000000
Rwpos68_78 in68_78 sp68_78 78000.000000
Rwpos68_79 in68_79 sp68_79 202000.000000
Rwpos68_80 in68_80 sp68_80 202000.000000
Rwpos68_81 in68_81 sp68_81 202000.000000
Rwpos68_82 in68_82 sp68_82 202000.000000
Rwpos68_83 in68_83 sp68_83 78000.000000
Rwpos68_84 in68_84 sp68_84 78000.000000
Rwpos69_1 in69_1 sp69_1 78000.000000
Rwpos69_2 in69_2 sp69_2 202000.000000
Rwpos69_3 in69_3 sp69_3 202000.000000
Rwpos69_4 in69_4 sp69_4 78000.000000
Rwpos69_5 in69_5 sp69_5 78000.000000
Rwpos69_6 in69_6 sp69_6 78000.000000
Rwpos69_7 in69_7 sp69_7 202000.000000
Rwpos69_8 in69_8 sp69_8 202000.000000
Rwpos69_9 in69_9 sp69_9 78000.000000
Rwpos69_10 in69_10 sp69_10 78000.000000
Rwpos69_11 in69_11 sp69_11 202000.000000
Rwpos69_12 in69_12 sp69_12 78000.000000
Rwpos69_13 in69_13 sp69_13 78000.000000
Rwpos69_14 in69_14 sp69_14 202000.000000
Rwpos69_15 in69_15 sp69_15 202000.000000
Rwpos69_16 in69_16 sp69_16 78000.000000
Rwpos69_17 in69_17 sp69_17 202000.000000
Rwpos69_18 in69_18 sp69_18 78000.000000
Rwpos69_19 in69_19 sp69_19 78000.000000
Rwpos69_20 in69_20 sp69_20 78000.000000
Rwpos69_21 in69_21 sp69_21 202000.000000
Rwpos69_22 in69_22 sp69_22 202000.000000
Rwpos69_23 in69_23 sp69_23 78000.000000
Rwpos69_24 in69_24 sp69_24 78000.000000
Rwpos69_25 in69_25 sp69_25 202000.000000
Rwpos69_26 in69_26 sp69_26 202000.000000
Rwpos69_27 in69_27 sp69_27 78000.000000
Rwpos69_28 in69_28 sp69_28 78000.000000
Rwpos69_29 in69_29 sp69_29 202000.000000
Rwpos69_30 in69_30 sp69_30 202000.000000
Rwpos69_31 in69_31 sp69_31 202000.000000
Rwpos69_32 in69_32 sp69_32 78000.000000
Rwpos69_33 in69_33 sp69_33 202000.000000
Rwpos69_34 in69_34 sp69_34 78000.000000
Rwpos69_35 in69_35 sp69_35 202000.000000
Rwpos69_36 in69_36 sp69_36 78000.000000
Rwpos69_37 in69_37 sp69_37 202000.000000
Rwpos69_38 in69_38 sp69_38 78000.000000
Rwpos69_39 in69_39 sp69_39 78000.000000
Rwpos69_40 in69_40 sp69_40 78000.000000
Rwpos69_41 in69_41 sp69_41 202000.000000
Rwpos69_42 in69_42 sp69_42 202000.000000
Rwpos69_43 in69_43 sp69_43 78000.000000
Rwpos69_44 in69_44 sp69_44 202000.000000
Rwpos69_45 in69_45 sp69_45 78000.000000
Rwpos69_46 in69_46 sp69_46 202000.000000
Rwpos69_47 in69_47 sp69_47 78000.000000
Rwpos69_48 in69_48 sp69_48 78000.000000
Rwpos69_49 in69_49 sp69_49 202000.000000
Rwpos69_50 in69_50 sp69_50 202000.000000
Rwpos69_51 in69_51 sp69_51 202000.000000
Rwpos69_52 in69_52 sp69_52 202000.000000
Rwpos69_53 in69_53 sp69_53 202000.000000
Rwpos69_54 in69_54 sp69_54 78000.000000
Rwpos69_55 in69_55 sp69_55 202000.000000
Rwpos69_56 in69_56 sp69_56 78000.000000
Rwpos69_57 in69_57 sp69_57 78000.000000
Rwpos69_58 in69_58 sp69_58 202000.000000
Rwpos69_59 in69_59 sp69_59 202000.000000
Rwpos69_60 in69_60 sp69_60 202000.000000
Rwpos69_61 in69_61 sp69_61 202000.000000
Rwpos69_62 in69_62 sp69_62 202000.000000
Rwpos69_63 in69_63 sp69_63 78000.000000
Rwpos69_64 in69_64 sp69_64 202000.000000
Rwpos69_65 in69_65 sp69_65 78000.000000
Rwpos69_66 in69_66 sp69_66 78000.000000
Rwpos69_67 in69_67 sp69_67 78000.000000
Rwpos69_68 in69_68 sp69_68 78000.000000
Rwpos69_69 in69_69 sp69_69 78000.000000
Rwpos69_70 in69_70 sp69_70 78000.000000
Rwpos69_71 in69_71 sp69_71 78000.000000
Rwpos69_72 in69_72 sp69_72 202000.000000
Rwpos69_73 in69_73 sp69_73 78000.000000
Rwpos69_74 in69_74 sp69_74 202000.000000
Rwpos69_75 in69_75 sp69_75 78000.000000
Rwpos69_76 in69_76 sp69_76 78000.000000
Rwpos69_77 in69_77 sp69_77 78000.000000
Rwpos69_78 in69_78 sp69_78 202000.000000
Rwpos69_79 in69_79 sp69_79 78000.000000
Rwpos69_80 in69_80 sp69_80 78000.000000
Rwpos69_81 in69_81 sp69_81 78000.000000
Rwpos69_82 in69_82 sp69_82 78000.000000
Rwpos69_83 in69_83 sp69_83 202000.000000
Rwpos69_84 in69_84 sp69_84 78000.000000
Rwpos70_1 in70_1 sp70_1 78000.000000
Rwpos70_2 in70_2 sp70_2 78000.000000
Rwpos70_3 in70_3 sp70_3 202000.000000
Rwpos70_4 in70_4 sp70_4 202000.000000
Rwpos70_5 in70_5 sp70_5 78000.000000
Rwpos70_6 in70_6 sp70_6 78000.000000
Rwpos70_7 in70_7 sp70_7 78000.000000
Rwpos70_8 in70_8 sp70_8 78000.000000
Rwpos70_9 in70_9 sp70_9 78000.000000
Rwpos70_10 in70_10 sp70_10 202000.000000
Rwpos70_11 in70_11 sp70_11 202000.000000
Rwpos70_12 in70_12 sp70_12 78000.000000
Rwpos70_13 in70_13 sp70_13 202000.000000
Rwpos70_14 in70_14 sp70_14 78000.000000
Rwpos70_15 in70_15 sp70_15 78000.000000
Rwpos70_16 in70_16 sp70_16 202000.000000
Rwpos70_17 in70_17 sp70_17 202000.000000
Rwpos70_18 in70_18 sp70_18 78000.000000
Rwpos70_19 in70_19 sp70_19 78000.000000
Rwpos70_20 in70_20 sp70_20 78000.000000
Rwpos70_21 in70_21 sp70_21 202000.000000
Rwpos70_22 in70_22 sp70_22 202000.000000
Rwpos70_23 in70_23 sp70_23 78000.000000
Rwpos70_24 in70_24 sp70_24 202000.000000
Rwpos70_25 in70_25 sp70_25 78000.000000
Rwpos70_26 in70_26 sp70_26 78000.000000
Rwpos70_27 in70_27 sp70_27 78000.000000
Rwpos70_28 in70_28 sp70_28 202000.000000
Rwpos70_29 in70_29 sp70_29 78000.000000
Rwpos70_30 in70_30 sp70_30 202000.000000
Rwpos70_31 in70_31 sp70_31 202000.000000
Rwpos70_32 in70_32 sp70_32 202000.000000
Rwpos70_33 in70_33 sp70_33 202000.000000
Rwpos70_34 in70_34 sp70_34 78000.000000
Rwpos70_35 in70_35 sp70_35 202000.000000
Rwpos70_36 in70_36 sp70_36 202000.000000
Rwpos70_37 in70_37 sp70_37 78000.000000
Rwpos70_38 in70_38 sp70_38 202000.000000
Rwpos70_39 in70_39 sp70_39 78000.000000
Rwpos70_40 in70_40 sp70_40 78000.000000
Rwpos70_41 in70_41 sp70_41 202000.000000
Rwpos70_42 in70_42 sp70_42 78000.000000
Rwpos70_43 in70_43 sp70_43 78000.000000
Rwpos70_44 in70_44 sp70_44 202000.000000
Rwpos70_45 in70_45 sp70_45 78000.000000
Rwpos70_46 in70_46 sp70_46 78000.000000
Rwpos70_47 in70_47 sp70_47 202000.000000
Rwpos70_48 in70_48 sp70_48 78000.000000
Rwpos70_49 in70_49 sp70_49 78000.000000
Rwpos70_50 in70_50 sp70_50 78000.000000
Rwpos70_51 in70_51 sp70_51 202000.000000
Rwpos70_52 in70_52 sp70_52 78000.000000
Rwpos70_53 in70_53 sp70_53 78000.000000
Rwpos70_54 in70_54 sp70_54 78000.000000
Rwpos70_55 in70_55 sp70_55 202000.000000
Rwpos70_56 in70_56 sp70_56 78000.000000
Rwpos70_57 in70_57 sp70_57 202000.000000
Rwpos70_58 in70_58 sp70_58 78000.000000
Rwpos70_59 in70_59 sp70_59 202000.000000
Rwpos70_60 in70_60 sp70_60 78000.000000
Rwpos70_61 in70_61 sp70_61 202000.000000
Rwpos70_62 in70_62 sp70_62 202000.000000
Rwpos70_63 in70_63 sp70_63 78000.000000
Rwpos70_64 in70_64 sp70_64 78000.000000
Rwpos70_65 in70_65 sp70_65 78000.000000
Rwpos70_66 in70_66 sp70_66 78000.000000
Rwpos70_67 in70_67 sp70_67 78000.000000
Rwpos70_68 in70_68 sp70_68 202000.000000
Rwpos70_69 in70_69 sp70_69 78000.000000
Rwpos70_70 in70_70 sp70_70 202000.000000
Rwpos70_71 in70_71 sp70_71 78000.000000
Rwpos70_72 in70_72 sp70_72 78000.000000
Rwpos70_73 in70_73 sp70_73 78000.000000
Rwpos70_74 in70_74 sp70_74 78000.000000
Rwpos70_75 in70_75 sp70_75 202000.000000
Rwpos70_76 in70_76 sp70_76 78000.000000
Rwpos70_77 in70_77 sp70_77 202000.000000
Rwpos70_78 in70_78 sp70_78 78000.000000
Rwpos70_79 in70_79 sp70_79 78000.000000
Rwpos70_80 in70_80 sp70_80 78000.000000
Rwpos70_81 in70_81 sp70_81 202000.000000
Rwpos70_82 in70_82 sp70_82 78000.000000
Rwpos70_83 in70_83 sp70_83 78000.000000
Rwpos70_84 in70_84 sp70_84 202000.000000
Rwpos71_1 in71_1 sp71_1 78000.000000
Rwpos71_2 in71_2 sp71_2 202000.000000
Rwpos71_3 in71_3 sp71_3 78000.000000
Rwpos71_4 in71_4 sp71_4 78000.000000
Rwpos71_5 in71_5 sp71_5 202000.000000
Rwpos71_6 in71_6 sp71_6 78000.000000
Rwpos71_7 in71_7 sp71_7 202000.000000
Rwpos71_8 in71_8 sp71_8 202000.000000
Rwpos71_9 in71_9 sp71_9 78000.000000
Rwpos71_10 in71_10 sp71_10 202000.000000
Rwpos71_11 in71_11 sp71_11 202000.000000
Rwpos71_12 in71_12 sp71_12 78000.000000
Rwpos71_13 in71_13 sp71_13 202000.000000
Rwpos71_14 in71_14 sp71_14 78000.000000
Rwpos71_15 in71_15 sp71_15 78000.000000
Rwpos71_16 in71_16 sp71_16 78000.000000
Rwpos71_17 in71_17 sp71_17 78000.000000
Rwpos71_18 in71_18 sp71_18 202000.000000
Rwpos71_19 in71_19 sp71_19 78000.000000
Rwpos71_20 in71_20 sp71_20 202000.000000
Rwpos71_21 in71_21 sp71_21 202000.000000
Rwpos71_22 in71_22 sp71_22 78000.000000
Rwpos71_23 in71_23 sp71_23 202000.000000
Rwpos71_24 in71_24 sp71_24 78000.000000
Rwpos71_25 in71_25 sp71_25 78000.000000
Rwpos71_26 in71_26 sp71_26 78000.000000
Rwpos71_27 in71_27 sp71_27 202000.000000
Rwpos71_28 in71_28 sp71_28 202000.000000
Rwpos71_29 in71_29 sp71_29 202000.000000
Rwpos71_30 in71_30 sp71_30 78000.000000
Rwpos71_31 in71_31 sp71_31 78000.000000
Rwpos71_32 in71_32 sp71_32 78000.000000
Rwpos71_33 in71_33 sp71_33 202000.000000
Rwpos71_34 in71_34 sp71_34 78000.000000
Rwpos71_35 in71_35 sp71_35 78000.000000
Rwpos71_36 in71_36 sp71_36 78000.000000
Rwpos71_37 in71_37 sp71_37 202000.000000
Rwpos71_38 in71_38 sp71_38 78000.000000
Rwpos71_39 in71_39 sp71_39 78000.000000
Rwpos71_40 in71_40 sp71_40 78000.000000
Rwpos71_41 in71_41 sp71_41 78000.000000
Rwpos71_42 in71_42 sp71_42 202000.000000
Rwpos71_43 in71_43 sp71_43 202000.000000
Rwpos71_44 in71_44 sp71_44 78000.000000
Rwpos71_45 in71_45 sp71_45 202000.000000
Rwpos71_46 in71_46 sp71_46 78000.000000
Rwpos71_47 in71_47 sp71_47 78000.000000
Rwpos71_48 in71_48 sp71_48 78000.000000
Rwpos71_49 in71_49 sp71_49 78000.000000
Rwpos71_50 in71_50 sp71_50 78000.000000
Rwpos71_51 in71_51 sp71_51 78000.000000
Rwpos71_52 in71_52 sp71_52 78000.000000
Rwpos71_53 in71_53 sp71_53 202000.000000
Rwpos71_54 in71_54 sp71_54 202000.000000
Rwpos71_55 in71_55 sp71_55 202000.000000
Rwpos71_56 in71_56 sp71_56 202000.000000
Rwpos71_57 in71_57 sp71_57 78000.000000
Rwpos71_58 in71_58 sp71_58 78000.000000
Rwpos71_59 in71_59 sp71_59 202000.000000
Rwpos71_60 in71_60 sp71_60 78000.000000
Rwpos71_61 in71_61 sp71_61 78000.000000
Rwpos71_62 in71_62 sp71_62 202000.000000
Rwpos71_63 in71_63 sp71_63 78000.000000
Rwpos71_64 in71_64 sp71_64 202000.000000
Rwpos71_65 in71_65 sp71_65 202000.000000
Rwpos71_66 in71_66 sp71_66 78000.000000
Rwpos71_67 in71_67 sp71_67 78000.000000
Rwpos71_68 in71_68 sp71_68 78000.000000
Rwpos71_69 in71_69 sp71_69 202000.000000
Rwpos71_70 in71_70 sp71_70 78000.000000
Rwpos71_71 in71_71 sp71_71 78000.000000
Rwpos71_72 in71_72 sp71_72 78000.000000
Rwpos71_73 in71_73 sp71_73 78000.000000
Rwpos71_74 in71_74 sp71_74 78000.000000
Rwpos71_75 in71_75 sp71_75 78000.000000
Rwpos71_76 in71_76 sp71_76 78000.000000
Rwpos71_77 in71_77 sp71_77 78000.000000
Rwpos71_78 in71_78 sp71_78 202000.000000
Rwpos71_79 in71_79 sp71_79 202000.000000
Rwpos71_80 in71_80 sp71_80 202000.000000
Rwpos71_81 in71_81 sp71_81 202000.000000
Rwpos71_82 in71_82 sp71_82 202000.000000
Rwpos71_83 in71_83 sp71_83 78000.000000
Rwpos71_84 in71_84 sp71_84 78000.000000
Rwpos72_1 in72_1 sp72_1 78000.000000
Rwpos72_2 in72_2 sp72_2 202000.000000
Rwpos72_3 in72_3 sp72_3 202000.000000
Rwpos72_4 in72_4 sp72_4 202000.000000
Rwpos72_5 in72_5 sp72_5 202000.000000
Rwpos72_6 in72_6 sp72_6 78000.000000
Rwpos72_7 in72_7 sp72_7 202000.000000
Rwpos72_8 in72_8 sp72_8 202000.000000
Rwpos72_9 in72_9 sp72_9 202000.000000
Rwpos72_10 in72_10 sp72_10 78000.000000
Rwpos72_11 in72_11 sp72_11 78000.000000
Rwpos72_12 in72_12 sp72_12 202000.000000
Rwpos72_13 in72_13 sp72_13 202000.000000
Rwpos72_14 in72_14 sp72_14 202000.000000
Rwpos72_15 in72_15 sp72_15 78000.000000
Rwpos72_16 in72_16 sp72_16 78000.000000
Rwpos72_17 in72_17 sp72_17 78000.000000
Rwpos72_18 in72_18 sp72_18 202000.000000
Rwpos72_19 in72_19 sp72_19 202000.000000
Rwpos72_20 in72_20 sp72_20 78000.000000
Rwpos72_21 in72_21 sp72_21 78000.000000
Rwpos72_22 in72_22 sp72_22 78000.000000
Rwpos72_23 in72_23 sp72_23 78000.000000
Rwpos72_24 in72_24 sp72_24 78000.000000
Rwpos72_25 in72_25 sp72_25 202000.000000
Rwpos72_26 in72_26 sp72_26 202000.000000
Rwpos72_27 in72_27 sp72_27 202000.000000
Rwpos72_28 in72_28 sp72_28 202000.000000
Rwpos72_29 in72_29 sp72_29 78000.000000
Rwpos72_30 in72_30 sp72_30 78000.000000
Rwpos72_31 in72_31 sp72_31 202000.000000
Rwpos72_32 in72_32 sp72_32 78000.000000
Rwpos72_33 in72_33 sp72_33 78000.000000
Rwpos72_34 in72_34 sp72_34 202000.000000
Rwpos72_35 in72_35 sp72_35 202000.000000
Rwpos72_36 in72_36 sp72_36 202000.000000
Rwpos72_37 in72_37 sp72_37 78000.000000
Rwpos72_38 in72_38 sp72_38 202000.000000
Rwpos72_39 in72_39 sp72_39 202000.000000
Rwpos72_40 in72_40 sp72_40 78000.000000
Rwpos72_41 in72_41 sp72_41 78000.000000
Rwpos72_42 in72_42 sp72_42 78000.000000
Rwpos72_43 in72_43 sp72_43 202000.000000
Rwpos72_44 in72_44 sp72_44 78000.000000
Rwpos72_45 in72_45 sp72_45 78000.000000
Rwpos72_46 in72_46 sp72_46 202000.000000
Rwpos72_47 in72_47 sp72_47 202000.000000
Rwpos72_48 in72_48 sp72_48 78000.000000
Rwpos72_49 in72_49 sp72_49 202000.000000
Rwpos72_50 in72_50 sp72_50 78000.000000
Rwpos72_51 in72_51 sp72_51 78000.000000
Rwpos72_52 in72_52 sp72_52 202000.000000
Rwpos72_53 in72_53 sp72_53 202000.000000
Rwpos72_54 in72_54 sp72_54 202000.000000
Rwpos72_55 in72_55 sp72_55 202000.000000
Rwpos72_56 in72_56 sp72_56 202000.000000
Rwpos72_57 in72_57 sp72_57 78000.000000
Rwpos72_58 in72_58 sp72_58 78000.000000
Rwpos72_59 in72_59 sp72_59 78000.000000
Rwpos72_60 in72_60 sp72_60 202000.000000
Rwpos72_61 in72_61 sp72_61 78000.000000
Rwpos72_62 in72_62 sp72_62 78000.000000
Rwpos72_63 in72_63 sp72_63 202000.000000
Rwpos72_64 in72_64 sp72_64 78000.000000
Rwpos72_65 in72_65 sp72_65 202000.000000
Rwpos72_66 in72_66 sp72_66 202000.000000
Rwpos72_67 in72_67 sp72_67 202000.000000
Rwpos72_68 in72_68 sp72_68 78000.000000
Rwpos72_69 in72_69 sp72_69 202000.000000
Rwpos72_70 in72_70 sp72_70 78000.000000
Rwpos72_71 in72_71 sp72_71 202000.000000
Rwpos72_72 in72_72 sp72_72 202000.000000
Rwpos72_73 in72_73 sp72_73 78000.000000
Rwpos72_74 in72_74 sp72_74 78000.000000
Rwpos72_75 in72_75 sp72_75 202000.000000
Rwpos72_76 in72_76 sp72_76 202000.000000
Rwpos72_77 in72_77 sp72_77 78000.000000
Rwpos72_78 in72_78 sp72_78 78000.000000
Rwpos72_79 in72_79 sp72_79 78000.000000
Rwpos72_80 in72_80 sp72_80 78000.000000
Rwpos72_81 in72_81 sp72_81 78000.000000
Rwpos72_82 in72_82 sp72_82 202000.000000
Rwpos72_83 in72_83 sp72_83 202000.000000
Rwpos72_84 in72_84 sp72_84 78000.000000
Rwpos73_1 in73_1 sp73_1 78000.000000
Rwpos73_2 in73_2 sp73_2 78000.000000
Rwpos73_3 in73_3 sp73_3 78000.000000
Rwpos73_4 in73_4 sp73_4 78000.000000
Rwpos73_5 in73_5 sp73_5 202000.000000
Rwpos73_6 in73_6 sp73_6 202000.000000
Rwpos73_7 in73_7 sp73_7 202000.000000
Rwpos73_8 in73_8 sp73_8 78000.000000
Rwpos73_9 in73_9 sp73_9 202000.000000
Rwpos73_10 in73_10 sp73_10 78000.000000
Rwpos73_11 in73_11 sp73_11 202000.000000
Rwpos73_12 in73_12 sp73_12 202000.000000
Rwpos73_13 in73_13 sp73_13 202000.000000
Rwpos73_14 in73_14 sp73_14 78000.000000
Rwpos73_15 in73_15 sp73_15 202000.000000
Rwpos73_16 in73_16 sp73_16 202000.000000
Rwpos73_17 in73_17 sp73_17 202000.000000
Rwpos73_18 in73_18 sp73_18 78000.000000
Rwpos73_19 in73_19 sp73_19 202000.000000
Rwpos73_20 in73_20 sp73_20 78000.000000
Rwpos73_21 in73_21 sp73_21 202000.000000
Rwpos73_22 in73_22 sp73_22 78000.000000
Rwpos73_23 in73_23 sp73_23 202000.000000
Rwpos73_24 in73_24 sp73_24 78000.000000
Rwpos73_25 in73_25 sp73_25 78000.000000
Rwpos73_26 in73_26 sp73_26 202000.000000
Rwpos73_27 in73_27 sp73_27 78000.000000
Rwpos73_28 in73_28 sp73_28 202000.000000
Rwpos73_29 in73_29 sp73_29 202000.000000
Rwpos73_30 in73_30 sp73_30 78000.000000
Rwpos73_31 in73_31 sp73_31 202000.000000
Rwpos73_32 in73_32 sp73_32 78000.000000
Rwpos73_33 in73_33 sp73_33 78000.000000
Rwpos73_34 in73_34 sp73_34 78000.000000
Rwpos73_35 in73_35 sp73_35 78000.000000
Rwpos73_36 in73_36 sp73_36 78000.000000
Rwpos73_37 in73_37 sp73_37 202000.000000
Rwpos73_38 in73_38 sp73_38 202000.000000
Rwpos73_39 in73_39 sp73_39 202000.000000
Rwpos73_40 in73_40 sp73_40 202000.000000
Rwpos73_41 in73_41 sp73_41 202000.000000
Rwpos73_42 in73_42 sp73_42 202000.000000
Rwpos73_43 in73_43 sp73_43 78000.000000
Rwpos73_44 in73_44 sp73_44 202000.000000
Rwpos73_45 in73_45 sp73_45 202000.000000
Rwpos73_46 in73_46 sp73_46 78000.000000
Rwpos73_47 in73_47 sp73_47 202000.000000
Rwpos73_48 in73_48 sp73_48 202000.000000
Rwpos73_49 in73_49 sp73_49 78000.000000
Rwpos73_50 in73_50 sp73_50 202000.000000
Rwpos73_51 in73_51 sp73_51 202000.000000
Rwpos73_52 in73_52 sp73_52 78000.000000
Rwpos73_53 in73_53 sp73_53 202000.000000
Rwpos73_54 in73_54 sp73_54 202000.000000
Rwpos73_55 in73_55 sp73_55 202000.000000
Rwpos73_56 in73_56 sp73_56 78000.000000
Rwpos73_57 in73_57 sp73_57 78000.000000
Rwpos73_58 in73_58 sp73_58 78000.000000
Rwpos73_59 in73_59 sp73_59 202000.000000
Rwpos73_60 in73_60 sp73_60 78000.000000
Rwpos73_61 in73_61 sp73_61 78000.000000
Rwpos73_62 in73_62 sp73_62 202000.000000
Rwpos73_63 in73_63 sp73_63 202000.000000
Rwpos73_64 in73_64 sp73_64 202000.000000
Rwpos73_65 in73_65 sp73_65 202000.000000
Rwpos73_66 in73_66 sp73_66 78000.000000
Rwpos73_67 in73_67 sp73_67 78000.000000
Rwpos73_68 in73_68 sp73_68 202000.000000
Rwpos73_69 in73_69 sp73_69 78000.000000
Rwpos73_70 in73_70 sp73_70 202000.000000
Rwpos73_71 in73_71 sp73_71 78000.000000
Rwpos73_72 in73_72 sp73_72 78000.000000
Rwpos73_73 in73_73 sp73_73 78000.000000
Rwpos73_74 in73_74 sp73_74 78000.000000
Rwpos73_75 in73_75 sp73_75 78000.000000
Rwpos73_76 in73_76 sp73_76 78000.000000
Rwpos73_77 in73_77 sp73_77 78000.000000
Rwpos73_78 in73_78 sp73_78 78000.000000
Rwpos73_79 in73_79 sp73_79 202000.000000
Rwpos73_80 in73_80 sp73_80 202000.000000
Rwpos73_81 in73_81 sp73_81 202000.000000
Rwpos73_82 in73_82 sp73_82 202000.000000
Rwpos73_83 in73_83 sp73_83 78000.000000
Rwpos73_84 in73_84 sp73_84 78000.000000
Rwpos74_1 in74_1 sp74_1 78000.000000
Rwpos74_2 in74_2 sp74_2 78000.000000
Rwpos74_3 in74_3 sp74_3 78000.000000
Rwpos74_4 in74_4 sp74_4 202000.000000
Rwpos74_5 in74_5 sp74_5 202000.000000
Rwpos74_6 in74_6 sp74_6 78000.000000
Rwpos74_7 in74_7 sp74_7 78000.000000
Rwpos74_8 in74_8 sp74_8 202000.000000
Rwpos74_9 in74_9 sp74_9 202000.000000
Rwpos74_10 in74_10 sp74_10 78000.000000
Rwpos74_11 in74_11 sp74_11 202000.000000
Rwpos74_12 in74_12 sp74_12 202000.000000
Rwpos74_13 in74_13 sp74_13 202000.000000
Rwpos74_14 in74_14 sp74_14 78000.000000
Rwpos74_15 in74_15 sp74_15 202000.000000
Rwpos74_16 in74_16 sp74_16 202000.000000
Rwpos74_17 in74_17 sp74_17 202000.000000
Rwpos74_18 in74_18 sp74_18 202000.000000
Rwpos74_19 in74_19 sp74_19 202000.000000
Rwpos74_20 in74_20 sp74_20 78000.000000
Rwpos74_21 in74_21 sp74_21 78000.000000
Rwpos74_22 in74_22 sp74_22 202000.000000
Rwpos74_23 in74_23 sp74_23 78000.000000
Rwpos74_24 in74_24 sp74_24 78000.000000
Rwpos74_25 in74_25 sp74_25 78000.000000
Rwpos74_26 in74_26 sp74_26 202000.000000
Rwpos74_27 in74_27 sp74_27 202000.000000
Rwpos74_28 in74_28 sp74_28 202000.000000
Rwpos74_29 in74_29 sp74_29 202000.000000
Rwpos74_30 in74_30 sp74_30 78000.000000
Rwpos74_31 in74_31 sp74_31 202000.000000
Rwpos74_32 in74_32 sp74_32 78000.000000
Rwpos74_33 in74_33 sp74_33 202000.000000
Rwpos74_34 in74_34 sp74_34 78000.000000
Rwpos74_35 in74_35 sp74_35 202000.000000
Rwpos74_36 in74_36 sp74_36 78000.000000
Rwpos74_37 in74_37 sp74_37 78000.000000
Rwpos74_38 in74_38 sp74_38 78000.000000
Rwpos74_39 in74_39 sp74_39 202000.000000
Rwpos74_40 in74_40 sp74_40 78000.000000
Rwpos74_41 in74_41 sp74_41 78000.000000
Rwpos74_42 in74_42 sp74_42 78000.000000
Rwpos74_43 in74_43 sp74_43 78000.000000
Rwpos74_44 in74_44 sp74_44 202000.000000
Rwpos74_45 in74_45 sp74_45 202000.000000
Rwpos74_46 in74_46 sp74_46 78000.000000
Rwpos74_47 in74_47 sp74_47 78000.000000
Rwpos74_48 in74_48 sp74_48 78000.000000
Rwpos74_49 in74_49 sp74_49 78000.000000
Rwpos74_50 in74_50 sp74_50 78000.000000
Rwpos74_51 in74_51 sp74_51 78000.000000
Rwpos74_52 in74_52 sp74_52 78000.000000
Rwpos74_53 in74_53 sp74_53 78000.000000
Rwpos74_54 in74_54 sp74_54 202000.000000
Rwpos74_55 in74_55 sp74_55 202000.000000
Rwpos74_56 in74_56 sp74_56 78000.000000
Rwpos74_57 in74_57 sp74_57 202000.000000
Rwpos74_58 in74_58 sp74_58 202000.000000
Rwpos74_59 in74_59 sp74_59 78000.000000
Rwpos74_60 in74_60 sp74_60 78000.000000
Rwpos74_61 in74_61 sp74_61 202000.000000
Rwpos74_62 in74_62 sp74_62 78000.000000
Rwpos74_63 in74_63 sp74_63 78000.000000
Rwpos74_64 in74_64 sp74_64 202000.000000
Rwpos74_65 in74_65 sp74_65 202000.000000
Rwpos74_66 in74_66 sp74_66 78000.000000
Rwpos74_67 in74_67 sp74_67 202000.000000
Rwpos74_68 in74_68 sp74_68 202000.000000
Rwpos74_69 in74_69 sp74_69 78000.000000
Rwpos74_70 in74_70 sp74_70 202000.000000
Rwpos74_71 in74_71 sp74_71 78000.000000
Rwpos74_72 in74_72 sp74_72 202000.000000
Rwpos74_73 in74_73 sp74_73 78000.000000
Rwpos74_74 in74_74 sp74_74 202000.000000
Rwpos74_75 in74_75 sp74_75 202000.000000
Rwpos74_76 in74_76 sp74_76 78000.000000
Rwpos74_77 in74_77 sp74_77 202000.000000
Rwpos74_78 in74_78 sp74_78 78000.000000
Rwpos74_79 in74_79 sp74_79 78000.000000
Rwpos74_80 in74_80 sp74_80 202000.000000
Rwpos74_81 in74_81 sp74_81 78000.000000
Rwpos74_82 in74_82 sp74_82 78000.000000
Rwpos74_83 in74_83 sp74_83 78000.000000
Rwpos74_84 in74_84 sp74_84 78000.000000
Rwpos75_1 in75_1 sp75_1 78000.000000
Rwpos75_2 in75_2 sp75_2 202000.000000
Rwpos75_3 in75_3 sp75_3 202000.000000
Rwpos75_4 in75_4 sp75_4 202000.000000
Rwpos75_5 in75_5 sp75_5 202000.000000
Rwpos75_6 in75_6 sp75_6 202000.000000
Rwpos75_7 in75_7 sp75_7 78000.000000
Rwpos75_8 in75_8 sp75_8 78000.000000
Rwpos75_9 in75_9 sp75_9 78000.000000
Rwpos75_10 in75_10 sp75_10 78000.000000
Rwpos75_11 in75_11 sp75_11 202000.000000
Rwpos75_12 in75_12 sp75_12 78000.000000
Rwpos75_13 in75_13 sp75_13 202000.000000
Rwpos75_14 in75_14 sp75_14 78000.000000
Rwpos75_15 in75_15 sp75_15 202000.000000
Rwpos75_16 in75_16 sp75_16 202000.000000
Rwpos75_17 in75_17 sp75_17 78000.000000
Rwpos75_18 in75_18 sp75_18 202000.000000
Rwpos75_19 in75_19 sp75_19 202000.000000
Rwpos75_20 in75_20 sp75_20 202000.000000
Rwpos75_21 in75_21 sp75_21 202000.000000
Rwpos75_22 in75_22 sp75_22 78000.000000
Rwpos75_23 in75_23 sp75_23 78000.000000
Rwpos75_24 in75_24 sp75_24 202000.000000
Rwpos75_25 in75_25 sp75_25 202000.000000
Rwpos75_26 in75_26 sp75_26 78000.000000
Rwpos75_27 in75_27 sp75_27 78000.000000
Rwpos75_28 in75_28 sp75_28 202000.000000
Rwpos75_29 in75_29 sp75_29 202000.000000
Rwpos75_30 in75_30 sp75_30 202000.000000
Rwpos75_31 in75_31 sp75_31 78000.000000
Rwpos75_32 in75_32 sp75_32 78000.000000
Rwpos75_33 in75_33 sp75_33 202000.000000
Rwpos75_34 in75_34 sp75_34 78000.000000
Rwpos75_35 in75_35 sp75_35 78000.000000
Rwpos75_36 in75_36 sp75_36 202000.000000
Rwpos75_37 in75_37 sp75_37 78000.000000
Rwpos75_38 in75_38 sp75_38 202000.000000
Rwpos75_39 in75_39 sp75_39 202000.000000
Rwpos75_40 in75_40 sp75_40 202000.000000
Rwpos75_41 in75_41 sp75_41 78000.000000
Rwpos75_42 in75_42 sp75_42 78000.000000
Rwpos75_43 in75_43 sp75_43 202000.000000
Rwpos75_44 in75_44 sp75_44 202000.000000
Rwpos75_45 in75_45 sp75_45 202000.000000
Rwpos75_46 in75_46 sp75_46 78000.000000
Rwpos75_47 in75_47 sp75_47 202000.000000
Rwpos75_48 in75_48 sp75_48 202000.000000
Rwpos75_49 in75_49 sp75_49 78000.000000
Rwpos75_50 in75_50 sp75_50 202000.000000
Rwpos75_51 in75_51 sp75_51 78000.000000
Rwpos75_52 in75_52 sp75_52 202000.000000
Rwpos75_53 in75_53 sp75_53 202000.000000
Rwpos75_54 in75_54 sp75_54 202000.000000
Rwpos75_55 in75_55 sp75_55 202000.000000
Rwpos75_56 in75_56 sp75_56 78000.000000
Rwpos75_57 in75_57 sp75_57 202000.000000
Rwpos75_58 in75_58 sp75_58 78000.000000
Rwpos75_59 in75_59 sp75_59 78000.000000
Rwpos75_60 in75_60 sp75_60 78000.000000
Rwpos75_61 in75_61 sp75_61 78000.000000
Rwpos75_62 in75_62 sp75_62 78000.000000
Rwpos75_63 in75_63 sp75_63 78000.000000
Rwpos75_64 in75_64 sp75_64 78000.000000
Rwpos75_65 in75_65 sp75_65 202000.000000
Rwpos75_66 in75_66 sp75_66 78000.000000
Rwpos75_67 in75_67 sp75_67 202000.000000
Rwpos75_68 in75_68 sp75_68 78000.000000
Rwpos75_69 in75_69 sp75_69 78000.000000
Rwpos75_70 in75_70 sp75_70 202000.000000
Rwpos75_71 in75_71 sp75_71 202000.000000
Rwpos75_72 in75_72 sp75_72 78000.000000
Rwpos75_73 in75_73 sp75_73 78000.000000
Rwpos75_74 in75_74 sp75_74 78000.000000
Rwpos75_75 in75_75 sp75_75 202000.000000
Rwpos75_76 in75_76 sp75_76 78000.000000
Rwpos75_77 in75_77 sp75_77 202000.000000
Rwpos75_78 in75_78 sp75_78 78000.000000
Rwpos75_79 in75_79 sp75_79 78000.000000
Rwpos75_80 in75_80 sp75_80 78000.000000
Rwpos75_81 in75_81 sp75_81 202000.000000
Rwpos75_82 in75_82 sp75_82 78000.000000
Rwpos75_83 in75_83 sp75_83 202000.000000
Rwpos75_84 in75_84 sp75_84 202000.000000
Rwpos76_1 in76_1 sp76_1 202000.000000
Rwpos76_2 in76_2 sp76_2 78000.000000
Rwpos76_3 in76_3 sp76_3 202000.000000
Rwpos76_4 in76_4 sp76_4 202000.000000
Rwpos76_5 in76_5 sp76_5 78000.000000
Rwpos76_6 in76_6 sp76_6 202000.000000
Rwpos76_7 in76_7 sp76_7 78000.000000
Rwpos76_8 in76_8 sp76_8 202000.000000
Rwpos76_9 in76_9 sp76_9 202000.000000
Rwpos76_10 in76_10 sp76_10 78000.000000
Rwpos76_11 in76_11 sp76_11 78000.000000
Rwpos76_12 in76_12 sp76_12 202000.000000
Rwpos76_13 in76_13 sp76_13 202000.000000
Rwpos76_14 in76_14 sp76_14 202000.000000
Rwpos76_15 in76_15 sp76_15 78000.000000
Rwpos76_16 in76_16 sp76_16 202000.000000
Rwpos76_17 in76_17 sp76_17 78000.000000
Rwpos76_18 in76_18 sp76_18 202000.000000
Rwpos76_19 in76_19 sp76_19 78000.000000
Rwpos76_20 in76_20 sp76_20 78000.000000
Rwpos76_21 in76_21 sp76_21 202000.000000
Rwpos76_22 in76_22 sp76_22 202000.000000
Rwpos76_23 in76_23 sp76_23 202000.000000
Rwpos76_24 in76_24 sp76_24 78000.000000
Rwpos76_25 in76_25 sp76_25 78000.000000
Rwpos76_26 in76_26 sp76_26 202000.000000
Rwpos76_27 in76_27 sp76_27 202000.000000
Rwpos76_28 in76_28 sp76_28 78000.000000
Rwpos76_29 in76_29 sp76_29 202000.000000
Rwpos76_30 in76_30 sp76_30 78000.000000
Rwpos76_31 in76_31 sp76_31 202000.000000
Rwpos76_32 in76_32 sp76_32 78000.000000
Rwpos76_33 in76_33 sp76_33 78000.000000
Rwpos76_34 in76_34 sp76_34 78000.000000
Rwpos76_35 in76_35 sp76_35 202000.000000
Rwpos76_36 in76_36 sp76_36 78000.000000
Rwpos76_37 in76_37 sp76_37 78000.000000
Rwpos76_38 in76_38 sp76_38 202000.000000
Rwpos76_39 in76_39 sp76_39 202000.000000
Rwpos76_40 in76_40 sp76_40 202000.000000
Rwpos76_41 in76_41 sp76_41 202000.000000
Rwpos76_42 in76_42 sp76_42 78000.000000
Rwpos76_43 in76_43 sp76_43 202000.000000
Rwpos76_44 in76_44 sp76_44 78000.000000
Rwpos76_45 in76_45 sp76_45 202000.000000
Rwpos76_46 in76_46 sp76_46 78000.000000
Rwpos76_47 in76_47 sp76_47 78000.000000
Rwpos76_48 in76_48 sp76_48 202000.000000
Rwpos76_49 in76_49 sp76_49 78000.000000
Rwpos76_50 in76_50 sp76_50 78000.000000
Rwpos76_51 in76_51 sp76_51 78000.000000
Rwpos76_52 in76_52 sp76_52 78000.000000
Rwpos76_53 in76_53 sp76_53 78000.000000
Rwpos76_54 in76_54 sp76_54 78000.000000
Rwpos76_55 in76_55 sp76_55 78000.000000
Rwpos76_56 in76_56 sp76_56 78000.000000
Rwpos76_57 in76_57 sp76_57 202000.000000
Rwpos76_58 in76_58 sp76_58 202000.000000
Rwpos76_59 in76_59 sp76_59 202000.000000
Rwpos76_60 in76_60 sp76_60 78000.000000
Rwpos76_61 in76_61 sp76_61 78000.000000
Rwpos76_62 in76_62 sp76_62 78000.000000
Rwpos76_63 in76_63 sp76_63 202000.000000
Rwpos76_64 in76_64 sp76_64 78000.000000
Rwpos76_65 in76_65 sp76_65 202000.000000
Rwpos76_66 in76_66 sp76_66 78000.000000
Rwpos76_67 in76_67 sp76_67 202000.000000
Rwpos76_68 in76_68 sp76_68 202000.000000
Rwpos76_69 in76_69 sp76_69 78000.000000
Rwpos76_70 in76_70 sp76_70 202000.000000
Rwpos76_71 in76_71 sp76_71 202000.000000
Rwpos76_72 in76_72 sp76_72 202000.000000
Rwpos76_73 in76_73 sp76_73 202000.000000
Rwpos76_74 in76_74 sp76_74 202000.000000
Rwpos76_75 in76_75 sp76_75 202000.000000
Rwpos76_76 in76_76 sp76_76 78000.000000
Rwpos76_77 in76_77 sp76_77 202000.000000
Rwpos76_78 in76_78 sp76_78 78000.000000
Rwpos76_79 in76_79 sp76_79 78000.000000
Rwpos76_80 in76_80 sp76_80 78000.000000
Rwpos76_81 in76_81 sp76_81 78000.000000
Rwpos76_82 in76_82 sp76_82 78000.000000
Rwpos76_83 in76_83 sp76_83 202000.000000
Rwpos76_84 in76_84 sp76_84 202000.000000
Rwpos77_1 in77_1 sp77_1 78000.000000
Rwpos77_2 in77_2 sp77_2 78000.000000
Rwpos77_3 in77_3 sp77_3 78000.000000
Rwpos77_4 in77_4 sp77_4 78000.000000
Rwpos77_5 in77_5 sp77_5 78000.000000
Rwpos77_6 in77_6 sp77_6 202000.000000
Rwpos77_7 in77_7 sp77_7 78000.000000
Rwpos77_8 in77_8 sp77_8 78000.000000
Rwpos77_9 in77_9 sp77_9 202000.000000
Rwpos77_10 in77_10 sp77_10 78000.000000
Rwpos77_11 in77_11 sp77_11 78000.000000
Rwpos77_12 in77_12 sp77_12 78000.000000
Rwpos77_13 in77_13 sp77_13 78000.000000
Rwpos77_14 in77_14 sp77_14 78000.000000
Rwpos77_15 in77_15 sp77_15 78000.000000
Rwpos77_16 in77_16 sp77_16 202000.000000
Rwpos77_17 in77_17 sp77_17 78000.000000
Rwpos77_18 in77_18 sp77_18 202000.000000
Rwpos77_19 in77_19 sp77_19 202000.000000
Rwpos77_20 in77_20 sp77_20 202000.000000
Rwpos77_21 in77_21 sp77_21 202000.000000
Rwpos77_22 in77_22 sp77_22 202000.000000
Rwpos77_23 in77_23 sp77_23 202000.000000
Rwpos77_24 in77_24 sp77_24 202000.000000
Rwpos77_25 in77_25 sp77_25 78000.000000
Rwpos77_26 in77_26 sp77_26 202000.000000
Rwpos77_27 in77_27 sp77_27 78000.000000
Rwpos77_28 in77_28 sp77_28 78000.000000
Rwpos77_29 in77_29 sp77_29 78000.000000
Rwpos77_30 in77_30 sp77_30 78000.000000
Rwpos77_31 in77_31 sp77_31 78000.000000
Rwpos77_32 in77_32 sp77_32 78000.000000
Rwpos77_33 in77_33 sp77_33 202000.000000
Rwpos77_34 in77_34 sp77_34 78000.000000
Rwpos77_35 in77_35 sp77_35 78000.000000
Rwpos77_36 in77_36 sp77_36 78000.000000
Rwpos77_37 in77_37 sp77_37 202000.000000
Rwpos77_38 in77_38 sp77_38 202000.000000
Rwpos77_39 in77_39 sp77_39 78000.000000
Rwpos77_40 in77_40 sp77_40 202000.000000
Rwpos77_41 in77_41 sp77_41 202000.000000
Rwpos77_42 in77_42 sp77_42 78000.000000
Rwpos77_43 in77_43 sp77_43 202000.000000
Rwpos77_44 in77_44 sp77_44 78000.000000
Rwpos77_45 in77_45 sp77_45 202000.000000
Rwpos77_46 in77_46 sp77_46 78000.000000
Rwpos77_47 in77_47 sp77_47 78000.000000
Rwpos77_48 in77_48 sp77_48 202000.000000
Rwpos77_49 in77_49 sp77_49 78000.000000
Rwpos77_50 in77_50 sp77_50 78000.000000
Rwpos77_51 in77_51 sp77_51 202000.000000
Rwpos77_52 in77_52 sp77_52 202000.000000
Rwpos77_53 in77_53 sp77_53 202000.000000
Rwpos77_54 in77_54 sp77_54 202000.000000
Rwpos77_55 in77_55 sp77_55 202000.000000
Rwpos77_56 in77_56 sp77_56 202000.000000
Rwpos77_57 in77_57 sp77_57 202000.000000
Rwpos77_58 in77_58 sp77_58 78000.000000
Rwpos77_59 in77_59 sp77_59 78000.000000
Rwpos77_60 in77_60 sp77_60 202000.000000
Rwpos77_61 in77_61 sp77_61 202000.000000
Rwpos77_62 in77_62 sp77_62 78000.000000
Rwpos77_63 in77_63 sp77_63 202000.000000
Rwpos77_64 in77_64 sp77_64 202000.000000
Rwpos77_65 in77_65 sp77_65 202000.000000
Rwpos77_66 in77_66 sp77_66 202000.000000
Rwpos77_67 in77_67 sp77_67 78000.000000
Rwpos77_68 in77_68 sp77_68 78000.000000
Rwpos77_69 in77_69 sp77_69 78000.000000
Rwpos77_70 in77_70 sp77_70 202000.000000
Rwpos77_71 in77_71 sp77_71 202000.000000
Rwpos77_72 in77_72 sp77_72 202000.000000
Rwpos77_73 in77_73 sp77_73 202000.000000
Rwpos77_74 in77_74 sp77_74 78000.000000
Rwpos77_75 in77_75 sp77_75 78000.000000
Rwpos77_76 in77_76 sp77_76 78000.000000
Rwpos77_77 in77_77 sp77_77 202000.000000
Rwpos77_78 in77_78 sp77_78 202000.000000
Rwpos77_79 in77_79 sp77_79 202000.000000
Rwpos77_80 in77_80 sp77_80 78000.000000
Rwpos77_81 in77_81 sp77_81 78000.000000
Rwpos77_82 in77_82 sp77_82 202000.000000
Rwpos77_83 in77_83 sp77_83 202000.000000
Rwpos77_84 in77_84 sp77_84 202000.000000
Rwpos78_1 in78_1 sp78_1 78000.000000
Rwpos78_2 in78_2 sp78_2 78000.000000
Rwpos78_3 in78_3 sp78_3 78000.000000
Rwpos78_4 in78_4 sp78_4 78000.000000
Rwpos78_5 in78_5 sp78_5 78000.000000
Rwpos78_6 in78_6 sp78_6 78000.000000
Rwpos78_7 in78_7 sp78_7 78000.000000
Rwpos78_8 in78_8 sp78_8 202000.000000
Rwpos78_9 in78_9 sp78_9 202000.000000
Rwpos78_10 in78_10 sp78_10 78000.000000
Rwpos78_11 in78_11 sp78_11 202000.000000
Rwpos78_12 in78_12 sp78_12 202000.000000
Rwpos78_13 in78_13 sp78_13 78000.000000
Rwpos78_14 in78_14 sp78_14 78000.000000
Rwpos78_15 in78_15 sp78_15 78000.000000
Rwpos78_16 in78_16 sp78_16 202000.000000
Rwpos78_17 in78_17 sp78_17 78000.000000
Rwpos78_18 in78_18 sp78_18 202000.000000
Rwpos78_19 in78_19 sp78_19 78000.000000
Rwpos78_20 in78_20 sp78_20 78000.000000
Rwpos78_21 in78_21 sp78_21 202000.000000
Rwpos78_22 in78_22 sp78_22 202000.000000
Rwpos78_23 in78_23 sp78_23 202000.000000
Rwpos78_24 in78_24 sp78_24 78000.000000
Rwpos78_25 in78_25 sp78_25 202000.000000
Rwpos78_26 in78_26 sp78_26 78000.000000
Rwpos78_27 in78_27 sp78_27 202000.000000
Rwpos78_28 in78_28 sp78_28 202000.000000
Rwpos78_29 in78_29 sp78_29 202000.000000
Rwpos78_30 in78_30 sp78_30 78000.000000
Rwpos78_31 in78_31 sp78_31 202000.000000
Rwpos78_32 in78_32 sp78_32 202000.000000
Rwpos78_33 in78_33 sp78_33 78000.000000
Rwpos78_34 in78_34 sp78_34 202000.000000
Rwpos78_35 in78_35 sp78_35 202000.000000
Rwpos78_36 in78_36 sp78_36 202000.000000
Rwpos78_37 in78_37 sp78_37 202000.000000
Rwpos78_38 in78_38 sp78_38 78000.000000
Rwpos78_39 in78_39 sp78_39 78000.000000
Rwpos78_40 in78_40 sp78_40 202000.000000
Rwpos78_41 in78_41 sp78_41 202000.000000
Rwpos78_42 in78_42 sp78_42 78000.000000
Rwpos78_43 in78_43 sp78_43 202000.000000
Rwpos78_44 in78_44 sp78_44 78000.000000
Rwpos78_45 in78_45 sp78_45 202000.000000
Rwpos78_46 in78_46 sp78_46 78000.000000
Rwpos78_47 in78_47 sp78_47 78000.000000
Rwpos78_48 in78_48 sp78_48 78000.000000
Rwpos78_49 in78_49 sp78_49 78000.000000
Rwpos78_50 in78_50 sp78_50 78000.000000
Rwpos78_51 in78_51 sp78_51 78000.000000
Rwpos78_52 in78_52 sp78_52 78000.000000
Rwpos78_53 in78_53 sp78_53 202000.000000
Rwpos78_54 in78_54 sp78_54 78000.000000
Rwpos78_55 in78_55 sp78_55 202000.000000
Rwpos78_56 in78_56 sp78_56 202000.000000
Rwpos78_57 in78_57 sp78_57 78000.000000
Rwpos78_58 in78_58 sp78_58 202000.000000
Rwpos78_59 in78_59 sp78_59 78000.000000
Rwpos78_60 in78_60 sp78_60 78000.000000
Rwpos78_61 in78_61 sp78_61 202000.000000
Rwpos78_62 in78_62 sp78_62 78000.000000
Rwpos78_63 in78_63 sp78_63 78000.000000
Rwpos78_64 in78_64 sp78_64 78000.000000
Rwpos78_65 in78_65 sp78_65 202000.000000
Rwpos78_66 in78_66 sp78_66 202000.000000
Rwpos78_67 in78_67 sp78_67 78000.000000
Rwpos78_68 in78_68 sp78_68 202000.000000
Rwpos78_69 in78_69 sp78_69 202000.000000
Rwpos78_70 in78_70 sp78_70 202000.000000
Rwpos78_71 in78_71 sp78_71 202000.000000
Rwpos78_72 in78_72 sp78_72 78000.000000
Rwpos78_73 in78_73 sp78_73 202000.000000
Rwpos78_74 in78_74 sp78_74 78000.000000
Rwpos78_75 in78_75 sp78_75 78000.000000
Rwpos78_76 in78_76 sp78_76 202000.000000
Rwpos78_77 in78_77 sp78_77 202000.000000
Rwpos78_78 in78_78 sp78_78 202000.000000
Rwpos78_79 in78_79 sp78_79 202000.000000
Rwpos78_80 in78_80 sp78_80 202000.000000
Rwpos78_81 in78_81 sp78_81 78000.000000
Rwpos78_82 in78_82 sp78_82 202000.000000
Rwpos78_83 in78_83 sp78_83 78000.000000
Rwpos78_84 in78_84 sp78_84 78000.000000
Rwpos79_1 in79_1 sp79_1 202000.000000
Rwpos79_2 in79_2 sp79_2 202000.000000
Rwpos79_3 in79_3 sp79_3 78000.000000
Rwpos79_4 in79_4 sp79_4 78000.000000
Rwpos79_5 in79_5 sp79_5 78000.000000
Rwpos79_6 in79_6 sp79_6 202000.000000
Rwpos79_7 in79_7 sp79_7 202000.000000
Rwpos79_8 in79_8 sp79_8 78000.000000
Rwpos79_9 in79_9 sp79_9 78000.000000
Rwpos79_10 in79_10 sp79_10 202000.000000
Rwpos79_11 in79_11 sp79_11 78000.000000
Rwpos79_12 in79_12 sp79_12 202000.000000
Rwpos79_13 in79_13 sp79_13 202000.000000
Rwpos79_14 in79_14 sp79_14 202000.000000
Rwpos79_15 in79_15 sp79_15 78000.000000
Rwpos79_16 in79_16 sp79_16 202000.000000
Rwpos79_17 in79_17 sp79_17 202000.000000
Rwpos79_18 in79_18 sp79_18 78000.000000
Rwpos79_19 in79_19 sp79_19 202000.000000
Rwpos79_20 in79_20 sp79_20 78000.000000
Rwpos79_21 in79_21 sp79_21 202000.000000
Rwpos79_22 in79_22 sp79_22 78000.000000
Rwpos79_23 in79_23 sp79_23 202000.000000
Rwpos79_24 in79_24 sp79_24 202000.000000
Rwpos79_25 in79_25 sp79_25 78000.000000
Rwpos79_26 in79_26 sp79_26 78000.000000
Rwpos79_27 in79_27 sp79_27 202000.000000
Rwpos79_28 in79_28 sp79_28 78000.000000
Rwpos79_29 in79_29 sp79_29 202000.000000
Rwpos79_30 in79_30 sp79_30 202000.000000
Rwpos79_31 in79_31 sp79_31 202000.000000
Rwpos79_32 in79_32 sp79_32 202000.000000
Rwpos79_33 in79_33 sp79_33 78000.000000
Rwpos79_34 in79_34 sp79_34 202000.000000
Rwpos79_35 in79_35 sp79_35 78000.000000
Rwpos79_36 in79_36 sp79_36 202000.000000
Rwpos79_37 in79_37 sp79_37 78000.000000
Rwpos79_38 in79_38 sp79_38 202000.000000
Rwpos79_39 in79_39 sp79_39 202000.000000
Rwpos79_40 in79_40 sp79_40 202000.000000
Rwpos79_41 in79_41 sp79_41 202000.000000
Rwpos79_42 in79_42 sp79_42 78000.000000
Rwpos79_43 in79_43 sp79_43 78000.000000
Rwpos79_44 in79_44 sp79_44 202000.000000
Rwpos79_45 in79_45 sp79_45 78000.000000
Rwpos79_46 in79_46 sp79_46 78000.000000
Rwpos79_47 in79_47 sp79_47 202000.000000
Rwpos79_48 in79_48 sp79_48 202000.000000
Rwpos79_49 in79_49 sp79_49 78000.000000
Rwpos79_50 in79_50 sp79_50 78000.000000
Rwpos79_51 in79_51 sp79_51 78000.000000
Rwpos79_52 in79_52 sp79_52 78000.000000
Rwpos79_53 in79_53 sp79_53 202000.000000
Rwpos79_54 in79_54 sp79_54 78000.000000
Rwpos79_55 in79_55 sp79_55 78000.000000
Rwpos79_56 in79_56 sp79_56 202000.000000
Rwpos79_57 in79_57 sp79_57 78000.000000
Rwpos79_58 in79_58 sp79_58 202000.000000
Rwpos79_59 in79_59 sp79_59 78000.000000
Rwpos79_60 in79_60 sp79_60 202000.000000
Rwpos79_61 in79_61 sp79_61 78000.000000
Rwpos79_62 in79_62 sp79_62 202000.000000
Rwpos79_63 in79_63 sp79_63 202000.000000
Rwpos79_64 in79_64 sp79_64 202000.000000
Rwpos79_65 in79_65 sp79_65 202000.000000
Rwpos79_66 in79_66 sp79_66 202000.000000
Rwpos79_67 in79_67 sp79_67 202000.000000
Rwpos79_68 in79_68 sp79_68 202000.000000
Rwpos79_69 in79_69 sp79_69 78000.000000
Rwpos79_70 in79_70 sp79_70 202000.000000
Rwpos79_71 in79_71 sp79_71 78000.000000
Rwpos79_72 in79_72 sp79_72 78000.000000
Rwpos79_73 in79_73 sp79_73 78000.000000
Rwpos79_74 in79_74 sp79_74 78000.000000
Rwpos79_75 in79_75 sp79_75 78000.000000
Rwpos79_76 in79_76 sp79_76 202000.000000
Rwpos79_77 in79_77 sp79_77 202000.000000
Rwpos79_78 in79_78 sp79_78 78000.000000
Rwpos79_79 in79_79 sp79_79 202000.000000
Rwpos79_80 in79_80 sp79_80 78000.000000
Rwpos79_81 in79_81 sp79_81 202000.000000
Rwpos79_82 in79_82 sp79_82 202000.000000
Rwpos79_83 in79_83 sp79_83 202000.000000
Rwpos79_84 in79_84 sp79_84 78000.000000
Rwpos80_1 in80_1 sp80_1 78000.000000
Rwpos80_2 in80_2 sp80_2 202000.000000
Rwpos80_3 in80_3 sp80_3 78000.000000
Rwpos80_4 in80_4 sp80_4 78000.000000
Rwpos80_5 in80_5 sp80_5 78000.000000
Rwpos80_6 in80_6 sp80_6 202000.000000
Rwpos80_7 in80_7 sp80_7 202000.000000
Rwpos80_8 in80_8 sp80_8 78000.000000
Rwpos80_9 in80_9 sp80_9 78000.000000
Rwpos80_10 in80_10 sp80_10 78000.000000
Rwpos80_11 in80_11 sp80_11 202000.000000
Rwpos80_12 in80_12 sp80_12 78000.000000
Rwpos80_13 in80_13 sp80_13 78000.000000
Rwpos80_14 in80_14 sp80_14 78000.000000
Rwpos80_15 in80_15 sp80_15 202000.000000
Rwpos80_16 in80_16 sp80_16 202000.000000
Rwpos80_17 in80_17 sp80_17 202000.000000
Rwpos80_18 in80_18 sp80_18 202000.000000
Rwpos80_19 in80_19 sp80_19 78000.000000
Rwpos80_20 in80_20 sp80_20 78000.000000
Rwpos80_21 in80_21 sp80_21 78000.000000
Rwpos80_22 in80_22 sp80_22 78000.000000
Rwpos80_23 in80_23 sp80_23 78000.000000
Rwpos80_24 in80_24 sp80_24 202000.000000
Rwpos80_25 in80_25 sp80_25 78000.000000
Rwpos80_26 in80_26 sp80_26 78000.000000
Rwpos80_27 in80_27 sp80_27 78000.000000
Rwpos80_28 in80_28 sp80_28 78000.000000
Rwpos80_29 in80_29 sp80_29 202000.000000
Rwpos80_30 in80_30 sp80_30 78000.000000
Rwpos80_31 in80_31 sp80_31 202000.000000
Rwpos80_32 in80_32 sp80_32 78000.000000
Rwpos80_33 in80_33 sp80_33 202000.000000
Rwpos80_34 in80_34 sp80_34 78000.000000
Rwpos80_35 in80_35 sp80_35 78000.000000
Rwpos80_36 in80_36 sp80_36 78000.000000
Rwpos80_37 in80_37 sp80_37 78000.000000
Rwpos80_38 in80_38 sp80_38 78000.000000
Rwpos80_39 in80_39 sp80_39 78000.000000
Rwpos80_40 in80_40 sp80_40 78000.000000
Rwpos80_41 in80_41 sp80_41 202000.000000
Rwpos80_42 in80_42 sp80_42 202000.000000
Rwpos80_43 in80_43 sp80_43 78000.000000
Rwpos80_44 in80_44 sp80_44 78000.000000
Rwpos80_45 in80_45 sp80_45 78000.000000
Rwpos80_46 in80_46 sp80_46 202000.000000
Rwpos80_47 in80_47 sp80_47 202000.000000
Rwpos80_48 in80_48 sp80_48 78000.000000
Rwpos80_49 in80_49 sp80_49 78000.000000
Rwpos80_50 in80_50 sp80_50 78000.000000
Rwpos80_51 in80_51 sp80_51 78000.000000
Rwpos80_52 in80_52 sp80_52 78000.000000
Rwpos80_53 in80_53 sp80_53 202000.000000
Rwpos80_54 in80_54 sp80_54 78000.000000
Rwpos80_55 in80_55 sp80_55 78000.000000
Rwpos80_56 in80_56 sp80_56 78000.000000
Rwpos80_57 in80_57 sp80_57 78000.000000
Rwpos80_58 in80_58 sp80_58 202000.000000
Rwpos80_59 in80_59 sp80_59 78000.000000
Rwpos80_60 in80_60 sp80_60 78000.000000
Rwpos80_61 in80_61 sp80_61 78000.000000
Rwpos80_62 in80_62 sp80_62 202000.000000
Rwpos80_63 in80_63 sp80_63 78000.000000
Rwpos80_64 in80_64 sp80_64 202000.000000
Rwpos80_65 in80_65 sp80_65 202000.000000
Rwpos80_66 in80_66 sp80_66 78000.000000
Rwpos80_67 in80_67 sp80_67 78000.000000
Rwpos80_68 in80_68 sp80_68 202000.000000
Rwpos80_69 in80_69 sp80_69 202000.000000
Rwpos80_70 in80_70 sp80_70 78000.000000
Rwpos80_71 in80_71 sp80_71 78000.000000
Rwpos80_72 in80_72 sp80_72 78000.000000
Rwpos80_73 in80_73 sp80_73 78000.000000
Rwpos80_74 in80_74 sp80_74 78000.000000
Rwpos80_75 in80_75 sp80_75 78000.000000
Rwpos80_76 in80_76 sp80_76 78000.000000
Rwpos80_77 in80_77 sp80_77 202000.000000
Rwpos80_78 in80_78 sp80_78 202000.000000
Rwpos80_79 in80_79 sp80_79 78000.000000
Rwpos80_80 in80_80 sp80_80 78000.000000
Rwpos80_81 in80_81 sp80_81 202000.000000
Rwpos80_82 in80_82 sp80_82 78000.000000
Rwpos80_83 in80_83 sp80_83 202000.000000
Rwpos80_84 in80_84 sp80_84 202000.000000
Rwpos81_1 in81_1 sp81_1 78000.000000
Rwpos81_2 in81_2 sp81_2 78000.000000
Rwpos81_3 in81_3 sp81_3 78000.000000
Rwpos81_4 in81_4 sp81_4 78000.000000
Rwpos81_5 in81_5 sp81_5 78000.000000
Rwpos81_6 in81_6 sp81_6 202000.000000
Rwpos81_7 in81_7 sp81_7 78000.000000
Rwpos81_8 in81_8 sp81_8 78000.000000
Rwpos81_9 in81_9 sp81_9 202000.000000
Rwpos81_10 in81_10 sp81_10 78000.000000
Rwpos81_11 in81_11 sp81_11 78000.000000
Rwpos81_12 in81_12 sp81_12 202000.000000
Rwpos81_13 in81_13 sp81_13 202000.000000
Rwpos81_14 in81_14 sp81_14 78000.000000
Rwpos81_15 in81_15 sp81_15 78000.000000
Rwpos81_16 in81_16 sp81_16 78000.000000
Rwpos81_17 in81_17 sp81_17 202000.000000
Rwpos81_18 in81_18 sp81_18 78000.000000
Rwpos81_19 in81_19 sp81_19 78000.000000
Rwpos81_20 in81_20 sp81_20 78000.000000
Rwpos81_21 in81_21 sp81_21 202000.000000
Rwpos81_22 in81_22 sp81_22 202000.000000
Rwpos81_23 in81_23 sp81_23 78000.000000
Rwpos81_24 in81_24 sp81_24 202000.000000
Rwpos81_25 in81_25 sp81_25 202000.000000
Rwpos81_26 in81_26 sp81_26 202000.000000
Rwpos81_27 in81_27 sp81_27 78000.000000
Rwpos81_28 in81_28 sp81_28 78000.000000
Rwpos81_29 in81_29 sp81_29 202000.000000
Rwpos81_30 in81_30 sp81_30 202000.000000
Rwpos81_31 in81_31 sp81_31 78000.000000
Rwpos81_32 in81_32 sp81_32 78000.000000
Rwpos81_33 in81_33 sp81_33 78000.000000
Rwpos81_34 in81_34 sp81_34 202000.000000
Rwpos81_35 in81_35 sp81_35 78000.000000
Rwpos81_36 in81_36 sp81_36 202000.000000
Rwpos81_37 in81_37 sp81_37 202000.000000
Rwpos81_38 in81_38 sp81_38 202000.000000
Rwpos81_39 in81_39 sp81_39 78000.000000
Rwpos81_40 in81_40 sp81_40 202000.000000
Rwpos81_41 in81_41 sp81_41 202000.000000
Rwpos81_42 in81_42 sp81_42 78000.000000
Rwpos81_43 in81_43 sp81_43 78000.000000
Rwpos81_44 in81_44 sp81_44 202000.000000
Rwpos81_45 in81_45 sp81_45 78000.000000
Rwpos81_46 in81_46 sp81_46 202000.000000
Rwpos81_47 in81_47 sp81_47 202000.000000
Rwpos81_48 in81_48 sp81_48 202000.000000
Rwpos81_49 in81_49 sp81_49 78000.000000
Rwpos81_50 in81_50 sp81_50 78000.000000
Rwpos81_51 in81_51 sp81_51 78000.000000
Rwpos81_52 in81_52 sp81_52 78000.000000
Rwpos81_53 in81_53 sp81_53 78000.000000
Rwpos81_54 in81_54 sp81_54 78000.000000
Rwpos81_55 in81_55 sp81_55 202000.000000
Rwpos81_56 in81_56 sp81_56 202000.000000
Rwpos81_57 in81_57 sp81_57 202000.000000
Rwpos81_58 in81_58 sp81_58 78000.000000
Rwpos81_59 in81_59 sp81_59 202000.000000
Rwpos81_60 in81_60 sp81_60 78000.000000
Rwpos81_61 in81_61 sp81_61 202000.000000
Rwpos81_62 in81_62 sp81_62 202000.000000
Rwpos81_63 in81_63 sp81_63 202000.000000
Rwpos81_64 in81_64 sp81_64 78000.000000
Rwpos81_65 in81_65 sp81_65 202000.000000
Rwpos81_66 in81_66 sp81_66 78000.000000
Rwpos81_67 in81_67 sp81_67 202000.000000
Rwpos81_68 in81_68 sp81_68 202000.000000
Rwpos81_69 in81_69 sp81_69 78000.000000
Rwpos81_70 in81_70 sp81_70 78000.000000
Rwpos81_71 in81_71 sp81_71 202000.000000
Rwpos81_72 in81_72 sp81_72 78000.000000
Rwpos81_73 in81_73 sp81_73 202000.000000
Rwpos81_74 in81_74 sp81_74 202000.000000
Rwpos81_75 in81_75 sp81_75 78000.000000
Rwpos81_76 in81_76 sp81_76 202000.000000
Rwpos81_77 in81_77 sp81_77 202000.000000
Rwpos81_78 in81_78 sp81_78 202000.000000
Rwpos81_79 in81_79 sp81_79 202000.000000
Rwpos81_80 in81_80 sp81_80 78000.000000
Rwpos81_81 in81_81 sp81_81 78000.000000
Rwpos81_82 in81_82 sp81_82 202000.000000
Rwpos81_83 in81_83 sp81_83 78000.000000
Rwpos81_84 in81_84 sp81_84 78000.000000
Rwpos82_1 in82_1 sp82_1 202000.000000
Rwpos82_2 in82_2 sp82_2 202000.000000
Rwpos82_3 in82_3 sp82_3 202000.000000
Rwpos82_4 in82_4 sp82_4 78000.000000
Rwpos82_5 in82_5 sp82_5 78000.000000
Rwpos82_6 in82_6 sp82_6 202000.000000
Rwpos82_7 in82_7 sp82_7 202000.000000
Rwpos82_8 in82_8 sp82_8 78000.000000
Rwpos82_9 in82_9 sp82_9 78000.000000
Rwpos82_10 in82_10 sp82_10 202000.000000
Rwpos82_11 in82_11 sp82_11 78000.000000
Rwpos82_12 in82_12 sp82_12 78000.000000
Rwpos82_13 in82_13 sp82_13 78000.000000
Rwpos82_14 in82_14 sp82_14 202000.000000
Rwpos82_15 in82_15 sp82_15 78000.000000
Rwpos82_16 in82_16 sp82_16 78000.000000
Rwpos82_17 in82_17 sp82_17 202000.000000
Rwpos82_18 in82_18 sp82_18 78000.000000
Rwpos82_19 in82_19 sp82_19 78000.000000
Rwpos82_20 in82_20 sp82_20 78000.000000
Rwpos82_21 in82_21 sp82_21 78000.000000
Rwpos82_22 in82_22 sp82_22 78000.000000
Rwpos82_23 in82_23 sp82_23 78000.000000
Rwpos82_24 in82_24 sp82_24 78000.000000
Rwpos82_25 in82_25 sp82_25 202000.000000
Rwpos82_26 in82_26 sp82_26 202000.000000
Rwpos82_27 in82_27 sp82_27 78000.000000
Rwpos82_28 in82_28 sp82_28 78000.000000
Rwpos82_29 in82_29 sp82_29 202000.000000
Rwpos82_30 in82_30 sp82_30 78000.000000
Rwpos82_31 in82_31 sp82_31 202000.000000
Rwpos82_32 in82_32 sp82_32 202000.000000
Rwpos82_33 in82_33 sp82_33 78000.000000
Rwpos82_34 in82_34 sp82_34 202000.000000
Rwpos82_35 in82_35 sp82_35 78000.000000
Rwpos82_36 in82_36 sp82_36 202000.000000
Rwpos82_37 in82_37 sp82_37 202000.000000
Rwpos82_38 in82_38 sp82_38 202000.000000
Rwpos82_39 in82_39 sp82_39 78000.000000
Rwpos82_40 in82_40 sp82_40 202000.000000
Rwpos82_41 in82_41 sp82_41 78000.000000
Rwpos82_42 in82_42 sp82_42 202000.000000
Rwpos82_43 in82_43 sp82_43 78000.000000
Rwpos82_44 in82_44 sp82_44 202000.000000
Rwpos82_45 in82_45 sp82_45 78000.000000
Rwpos82_46 in82_46 sp82_46 202000.000000
Rwpos82_47 in82_47 sp82_47 202000.000000
Rwpos82_48 in82_48 sp82_48 78000.000000
Rwpos82_49 in82_49 sp82_49 78000.000000
Rwpos82_50 in82_50 sp82_50 202000.000000
Rwpos82_51 in82_51 sp82_51 78000.000000
Rwpos82_52 in82_52 sp82_52 202000.000000
Rwpos82_53 in82_53 sp82_53 202000.000000
Rwpos82_54 in82_54 sp82_54 202000.000000
Rwpos82_55 in82_55 sp82_55 78000.000000
Rwpos82_56 in82_56 sp82_56 78000.000000
Rwpos82_57 in82_57 sp82_57 78000.000000
Rwpos82_58 in82_58 sp82_58 202000.000000
Rwpos82_59 in82_59 sp82_59 202000.000000
Rwpos82_60 in82_60 sp82_60 202000.000000
Rwpos82_61 in82_61 sp82_61 78000.000000
Rwpos82_62 in82_62 sp82_62 78000.000000
Rwpos82_63 in82_63 sp82_63 78000.000000
Rwpos82_64 in82_64 sp82_64 202000.000000
Rwpos82_65 in82_65 sp82_65 78000.000000
Rwpos82_66 in82_66 sp82_66 78000.000000
Rwpos82_67 in82_67 sp82_67 202000.000000
Rwpos82_68 in82_68 sp82_68 78000.000000
Rwpos82_69 in82_69 sp82_69 78000.000000
Rwpos82_70 in82_70 sp82_70 78000.000000
Rwpos82_71 in82_71 sp82_71 78000.000000
Rwpos82_72 in82_72 sp82_72 202000.000000
Rwpos82_73 in82_73 sp82_73 78000.000000
Rwpos82_74 in82_74 sp82_74 202000.000000
Rwpos82_75 in82_75 sp82_75 202000.000000
Rwpos82_76 in82_76 sp82_76 202000.000000
Rwpos82_77 in82_77 sp82_77 202000.000000
Rwpos82_78 in82_78 sp82_78 202000.000000
Rwpos82_79 in82_79 sp82_79 202000.000000
Rwpos82_80 in82_80 sp82_80 78000.000000
Rwpos82_81 in82_81 sp82_81 78000.000000
Rwpos82_82 in82_82 sp82_82 78000.000000
Rwpos82_83 in82_83 sp82_83 78000.000000
Rwpos82_84 in82_84 sp82_84 78000.000000
Rwpos83_1 in83_1 sp83_1 78000.000000
Rwpos83_2 in83_2 sp83_2 78000.000000
Rwpos83_3 in83_3 sp83_3 202000.000000
Rwpos83_4 in83_4 sp83_4 78000.000000
Rwpos83_5 in83_5 sp83_5 78000.000000
Rwpos83_6 in83_6 sp83_6 202000.000000
Rwpos83_7 in83_7 sp83_7 78000.000000
Rwpos83_8 in83_8 sp83_8 78000.000000
Rwpos83_9 in83_9 sp83_9 78000.000000
Rwpos83_10 in83_10 sp83_10 202000.000000
Rwpos83_11 in83_11 sp83_11 202000.000000
Rwpos83_12 in83_12 sp83_12 78000.000000
Rwpos83_13 in83_13 sp83_13 202000.000000
Rwpos83_14 in83_14 sp83_14 202000.000000
Rwpos83_15 in83_15 sp83_15 202000.000000
Rwpos83_16 in83_16 sp83_16 78000.000000
Rwpos83_17 in83_17 sp83_17 78000.000000
Rwpos83_18 in83_18 sp83_18 78000.000000
Rwpos83_19 in83_19 sp83_19 78000.000000
Rwpos83_20 in83_20 sp83_20 78000.000000
Rwpos83_21 in83_21 sp83_21 78000.000000
Rwpos83_22 in83_22 sp83_22 78000.000000
Rwpos83_23 in83_23 sp83_23 202000.000000
Rwpos83_24 in83_24 sp83_24 78000.000000
Rwpos83_25 in83_25 sp83_25 78000.000000
Rwpos83_26 in83_26 sp83_26 78000.000000
Rwpos83_27 in83_27 sp83_27 78000.000000
Rwpos83_28 in83_28 sp83_28 202000.000000
Rwpos83_29 in83_29 sp83_29 202000.000000
Rwpos83_30 in83_30 sp83_30 202000.000000
Rwpos83_31 in83_31 sp83_31 202000.000000
Rwpos83_32 in83_32 sp83_32 78000.000000
Rwpos83_33 in83_33 sp83_33 78000.000000
Rwpos83_34 in83_34 sp83_34 202000.000000
Rwpos83_35 in83_35 sp83_35 202000.000000
Rwpos83_36 in83_36 sp83_36 202000.000000
Rwpos83_37 in83_37 sp83_37 78000.000000
Rwpos83_38 in83_38 sp83_38 202000.000000
Rwpos83_39 in83_39 sp83_39 202000.000000
Rwpos83_40 in83_40 sp83_40 202000.000000
Rwpos83_41 in83_41 sp83_41 202000.000000
Rwpos83_42 in83_42 sp83_42 78000.000000
Rwpos83_43 in83_43 sp83_43 78000.000000
Rwpos83_44 in83_44 sp83_44 78000.000000
Rwpos83_45 in83_45 sp83_45 202000.000000
Rwpos83_46 in83_46 sp83_46 202000.000000
Rwpos83_47 in83_47 sp83_47 202000.000000
Rwpos83_48 in83_48 sp83_48 78000.000000
Rwpos83_49 in83_49 sp83_49 202000.000000
Rwpos83_50 in83_50 sp83_50 202000.000000
Rwpos83_51 in83_51 sp83_51 202000.000000
Rwpos83_52 in83_52 sp83_52 78000.000000
Rwpos83_53 in83_53 sp83_53 202000.000000
Rwpos83_54 in83_54 sp83_54 78000.000000
Rwpos83_55 in83_55 sp83_55 202000.000000
Rwpos83_56 in83_56 sp83_56 202000.000000
Rwpos83_57 in83_57 sp83_57 202000.000000
Rwpos83_58 in83_58 sp83_58 202000.000000
Rwpos83_59 in83_59 sp83_59 78000.000000
Rwpos83_60 in83_60 sp83_60 78000.000000
Rwpos83_61 in83_61 sp83_61 202000.000000
Rwpos83_62 in83_62 sp83_62 78000.000000
Rwpos83_63 in83_63 sp83_63 78000.000000
Rwpos83_64 in83_64 sp83_64 78000.000000
Rwpos83_65 in83_65 sp83_65 78000.000000
Rwpos83_66 in83_66 sp83_66 78000.000000
Rwpos83_67 in83_67 sp83_67 202000.000000
Rwpos83_68 in83_68 sp83_68 202000.000000
Rwpos83_69 in83_69 sp83_69 78000.000000
Rwpos83_70 in83_70 sp83_70 202000.000000
Rwpos83_71 in83_71 sp83_71 202000.000000
Rwpos83_72 in83_72 sp83_72 202000.000000
Rwpos83_73 in83_73 sp83_73 202000.000000
Rwpos83_74 in83_74 sp83_74 202000.000000
Rwpos83_75 in83_75 sp83_75 202000.000000
Rwpos83_76 in83_76 sp83_76 202000.000000
Rwpos83_77 in83_77 sp83_77 202000.000000
Rwpos83_78 in83_78 sp83_78 202000.000000
Rwpos83_79 in83_79 sp83_79 202000.000000
Rwpos83_80 in83_80 sp83_80 78000.000000
Rwpos83_81 in83_81 sp83_81 78000.000000
Rwpos83_82 in83_82 sp83_82 78000.000000
Rwpos83_83 in83_83 sp83_83 78000.000000
Rwpos83_84 in83_84 sp83_84 78000.000000
Rwpos84_1 in84_1 sp84_1 202000.000000
Rwpos84_2 in84_2 sp84_2 202000.000000
Rwpos84_3 in84_3 sp84_3 202000.000000
Rwpos84_4 in84_4 sp84_4 202000.000000
Rwpos84_5 in84_5 sp84_5 202000.000000
Rwpos84_6 in84_6 sp84_6 202000.000000
Rwpos84_7 in84_7 sp84_7 202000.000000
Rwpos84_8 in84_8 sp84_8 78000.000000
Rwpos84_9 in84_9 sp84_9 78000.000000
Rwpos84_10 in84_10 sp84_10 202000.000000
Rwpos84_11 in84_11 sp84_11 78000.000000
Rwpos84_12 in84_12 sp84_12 78000.000000
Rwpos84_13 in84_13 sp84_13 202000.000000
Rwpos84_14 in84_14 sp84_14 202000.000000
Rwpos84_15 in84_15 sp84_15 202000.000000
Rwpos84_16 in84_16 sp84_16 78000.000000
Rwpos84_17 in84_17 sp84_17 78000.000000
Rwpos84_18 in84_18 sp84_18 78000.000000
Rwpos84_19 in84_19 sp84_19 202000.000000
Rwpos84_20 in84_20 sp84_20 202000.000000
Rwpos84_21 in84_21 sp84_21 78000.000000
Rwpos84_22 in84_22 sp84_22 78000.000000
Rwpos84_23 in84_23 sp84_23 78000.000000
Rwpos84_24 in84_24 sp84_24 78000.000000
Rwpos84_25 in84_25 sp84_25 202000.000000
Rwpos84_26 in84_26 sp84_26 78000.000000
Rwpos84_27 in84_27 sp84_27 78000.000000
Rwpos84_28 in84_28 sp84_28 78000.000000
Rwpos84_29 in84_29 sp84_29 202000.000000
Rwpos84_30 in84_30 sp84_30 78000.000000
Rwpos84_31 in84_31 sp84_31 78000.000000
Rwpos84_32 in84_32 sp84_32 78000.000000
Rwpos84_33 in84_33 sp84_33 202000.000000
Rwpos84_34 in84_34 sp84_34 78000.000000
Rwpos84_35 in84_35 sp84_35 202000.000000
Rwpos84_36 in84_36 sp84_36 78000.000000
Rwpos84_37 in84_37 sp84_37 78000.000000
Rwpos84_38 in84_38 sp84_38 202000.000000
Rwpos84_39 in84_39 sp84_39 202000.000000
Rwpos84_40 in84_40 sp84_40 78000.000000
Rwpos84_41 in84_41 sp84_41 78000.000000
Rwpos84_42 in84_42 sp84_42 202000.000000
Rwpos84_43 in84_43 sp84_43 78000.000000
Rwpos84_44 in84_44 sp84_44 202000.000000
Rwpos84_45 in84_45 sp84_45 202000.000000
Rwpos84_46 in84_46 sp84_46 202000.000000
Rwpos84_47 in84_47 sp84_47 202000.000000
Rwpos84_48 in84_48 sp84_48 78000.000000
Rwpos84_49 in84_49 sp84_49 202000.000000
Rwpos84_50 in84_50 sp84_50 202000.000000
Rwpos84_51 in84_51 sp84_51 78000.000000
Rwpos84_52 in84_52 sp84_52 78000.000000
Rwpos84_53 in84_53 sp84_53 78000.000000
Rwpos84_54 in84_54 sp84_54 78000.000000
Rwpos84_55 in84_55 sp84_55 202000.000000
Rwpos84_56 in84_56 sp84_56 78000.000000
Rwpos84_57 in84_57 sp84_57 78000.000000
Rwpos84_58 in84_58 sp84_58 78000.000000
Rwpos84_59 in84_59 sp84_59 202000.000000
Rwpos84_60 in84_60 sp84_60 202000.000000
Rwpos84_61 in84_61 sp84_61 78000.000000
Rwpos84_62 in84_62 sp84_62 202000.000000
Rwpos84_63 in84_63 sp84_63 202000.000000
Rwpos84_64 in84_64 sp84_64 78000.000000
Rwpos84_65 in84_65 sp84_65 78000.000000
Rwpos84_66 in84_66 sp84_66 78000.000000
Rwpos84_67 in84_67 sp84_67 78000.000000
Rwpos84_68 in84_68 sp84_68 78000.000000
Rwpos84_69 in84_69 sp84_69 78000.000000
Rwpos84_70 in84_70 sp84_70 202000.000000
Rwpos84_71 in84_71 sp84_71 78000.000000
Rwpos84_72 in84_72 sp84_72 202000.000000
Rwpos84_73 in84_73 sp84_73 78000.000000
Rwpos84_74 in84_74 sp84_74 78000.000000
Rwpos84_75 in84_75 sp84_75 202000.000000
Rwpos84_76 in84_76 sp84_76 78000.000000
Rwpos84_77 in84_77 sp84_77 202000.000000
Rwpos84_78 in84_78 sp84_78 78000.000000
Rwpos84_79 in84_79 sp84_79 78000.000000
Rwpos84_80 in84_80 sp84_80 78000.000000
Rwpos84_81 in84_81 sp84_81 202000.000000
Rwpos84_82 in84_82 sp84_82 78000.000000
Rwpos84_83 in84_83 sp84_83 202000.000000
Rwpos84_84 in84_84 sp84_84 202000.000000
Rwpos85_1 in85_1 sp85_1 202000.000000
Rwpos85_2 in85_2 sp85_2 202000.000000
Rwpos85_3 in85_3 sp85_3 202000.000000
Rwpos85_4 in85_4 sp85_4 78000.000000
Rwpos85_5 in85_5 sp85_5 78000.000000
Rwpos85_6 in85_6 sp85_6 78000.000000
Rwpos85_7 in85_7 sp85_7 202000.000000
Rwpos85_8 in85_8 sp85_8 78000.000000
Rwpos85_9 in85_9 sp85_9 202000.000000
Rwpos85_10 in85_10 sp85_10 78000.000000
Rwpos85_11 in85_11 sp85_11 78000.000000
Rwpos85_12 in85_12 sp85_12 78000.000000
Rwpos85_13 in85_13 sp85_13 78000.000000
Rwpos85_14 in85_14 sp85_14 202000.000000
Rwpos85_15 in85_15 sp85_15 78000.000000
Rwpos85_16 in85_16 sp85_16 202000.000000
Rwpos85_17 in85_17 sp85_17 202000.000000
Rwpos85_18 in85_18 sp85_18 78000.000000
Rwpos85_19 in85_19 sp85_19 78000.000000
Rwpos85_20 in85_20 sp85_20 78000.000000
Rwpos85_21 in85_21 sp85_21 78000.000000
Rwpos85_22 in85_22 sp85_22 78000.000000
Rwpos85_23 in85_23 sp85_23 78000.000000
Rwpos85_24 in85_24 sp85_24 202000.000000
Rwpos85_25 in85_25 sp85_25 78000.000000
Rwpos85_26 in85_26 sp85_26 78000.000000
Rwpos85_27 in85_27 sp85_27 78000.000000
Rwpos85_28 in85_28 sp85_28 78000.000000
Rwpos85_29 in85_29 sp85_29 202000.000000
Rwpos85_30 in85_30 sp85_30 202000.000000
Rwpos85_31 in85_31 sp85_31 78000.000000
Rwpos85_32 in85_32 sp85_32 202000.000000
Rwpos85_33 in85_33 sp85_33 202000.000000
Rwpos85_34 in85_34 sp85_34 78000.000000
Rwpos85_35 in85_35 sp85_35 78000.000000
Rwpos85_36 in85_36 sp85_36 78000.000000
Rwpos85_37 in85_37 sp85_37 202000.000000
Rwpos85_38 in85_38 sp85_38 78000.000000
Rwpos85_39 in85_39 sp85_39 78000.000000
Rwpos85_40 in85_40 sp85_40 78000.000000
Rwpos85_41 in85_41 sp85_41 202000.000000
Rwpos85_42 in85_42 sp85_42 202000.000000
Rwpos85_43 in85_43 sp85_43 78000.000000
Rwpos85_44 in85_44 sp85_44 202000.000000
Rwpos85_45 in85_45 sp85_45 78000.000000
Rwpos85_46 in85_46 sp85_46 202000.000000
Rwpos85_47 in85_47 sp85_47 78000.000000
Rwpos85_48 in85_48 sp85_48 202000.000000
Rwpos85_49 in85_49 sp85_49 202000.000000
Rwpos85_50 in85_50 sp85_50 78000.000000
Rwpos85_51 in85_51 sp85_51 78000.000000
Rwpos85_52 in85_52 sp85_52 202000.000000
Rwpos85_53 in85_53 sp85_53 78000.000000
Rwpos85_54 in85_54 sp85_54 78000.000000
Rwpos85_55 in85_55 sp85_55 202000.000000
Rwpos85_56 in85_56 sp85_56 78000.000000
Rwpos85_57 in85_57 sp85_57 202000.000000
Rwpos85_58 in85_58 sp85_58 78000.000000
Rwpos85_59 in85_59 sp85_59 202000.000000
Rwpos85_60 in85_60 sp85_60 202000.000000
Rwpos85_61 in85_61 sp85_61 202000.000000
Rwpos85_62 in85_62 sp85_62 78000.000000
Rwpos85_63 in85_63 sp85_63 78000.000000
Rwpos85_64 in85_64 sp85_64 202000.000000
Rwpos85_65 in85_65 sp85_65 202000.000000
Rwpos85_66 in85_66 sp85_66 202000.000000
Rwpos85_67 in85_67 sp85_67 202000.000000
Rwpos85_68 in85_68 sp85_68 202000.000000
Rwpos85_69 in85_69 sp85_69 78000.000000
Rwpos85_70 in85_70 sp85_70 78000.000000
Rwpos85_71 in85_71 sp85_71 78000.000000
Rwpos85_72 in85_72 sp85_72 78000.000000
Rwpos85_73 in85_73 sp85_73 202000.000000
Rwpos85_74 in85_74 sp85_74 202000.000000
Rwpos85_75 in85_75 sp85_75 78000.000000
Rwpos85_76 in85_76 sp85_76 202000.000000
Rwpos85_77 in85_77 sp85_77 78000.000000
Rwpos85_78 in85_78 sp85_78 78000.000000
Rwpos85_79 in85_79 sp85_79 78000.000000
Rwpos85_80 in85_80 sp85_80 78000.000000
Rwpos85_81 in85_81 sp85_81 202000.000000
Rwpos85_82 in85_82 sp85_82 78000.000000
Rwpos85_83 in85_83 sp85_83 202000.000000
Rwpos85_84 in85_84 sp85_84 78000.000000
Rwpos86_1 in86_1 sp86_1 202000.000000
Rwpos86_2 in86_2 sp86_2 78000.000000
Rwpos86_3 in86_3 sp86_3 202000.000000
Rwpos86_4 in86_4 sp86_4 202000.000000
Rwpos86_5 in86_5 sp86_5 202000.000000
Rwpos86_6 in86_6 sp86_6 78000.000000
Rwpos86_7 in86_7 sp86_7 78000.000000
Rwpos86_8 in86_8 sp86_8 202000.000000
Rwpos86_9 in86_9 sp86_9 202000.000000
Rwpos86_10 in86_10 sp86_10 78000.000000
Rwpos86_11 in86_11 sp86_11 202000.000000
Rwpos86_12 in86_12 sp86_12 78000.000000
Rwpos86_13 in86_13 sp86_13 78000.000000
Rwpos86_14 in86_14 sp86_14 78000.000000
Rwpos86_15 in86_15 sp86_15 78000.000000
Rwpos86_16 in86_16 sp86_16 78000.000000
Rwpos86_17 in86_17 sp86_17 78000.000000
Rwpos86_18 in86_18 sp86_18 202000.000000
Rwpos86_19 in86_19 sp86_19 78000.000000
Rwpos86_20 in86_20 sp86_20 202000.000000
Rwpos86_21 in86_21 sp86_21 202000.000000
Rwpos86_22 in86_22 sp86_22 202000.000000
Rwpos86_23 in86_23 sp86_23 202000.000000
Rwpos86_24 in86_24 sp86_24 202000.000000
Rwpos86_25 in86_25 sp86_25 78000.000000
Rwpos86_26 in86_26 sp86_26 202000.000000
Rwpos86_27 in86_27 sp86_27 202000.000000
Rwpos86_28 in86_28 sp86_28 78000.000000
Rwpos86_29 in86_29 sp86_29 202000.000000
Rwpos86_30 in86_30 sp86_30 78000.000000
Rwpos86_31 in86_31 sp86_31 202000.000000
Rwpos86_32 in86_32 sp86_32 78000.000000
Rwpos86_33 in86_33 sp86_33 202000.000000
Rwpos86_34 in86_34 sp86_34 78000.000000
Rwpos86_35 in86_35 sp86_35 202000.000000
Rwpos86_36 in86_36 sp86_36 78000.000000
Rwpos86_37 in86_37 sp86_37 78000.000000
Rwpos86_38 in86_38 sp86_38 78000.000000
Rwpos86_39 in86_39 sp86_39 202000.000000
Rwpos86_40 in86_40 sp86_40 78000.000000
Rwpos86_41 in86_41 sp86_41 202000.000000
Rwpos86_42 in86_42 sp86_42 202000.000000
Rwpos86_43 in86_43 sp86_43 202000.000000
Rwpos86_44 in86_44 sp86_44 78000.000000
Rwpos86_45 in86_45 sp86_45 202000.000000
Rwpos86_46 in86_46 sp86_46 78000.000000
Rwpos86_47 in86_47 sp86_47 78000.000000
Rwpos86_48 in86_48 sp86_48 202000.000000
Rwpos86_49 in86_49 sp86_49 78000.000000
Rwpos86_50 in86_50 sp86_50 78000.000000
Rwpos86_51 in86_51 sp86_51 202000.000000
Rwpos86_52 in86_52 sp86_52 78000.000000
Rwpos86_53 in86_53 sp86_53 202000.000000
Rwpos86_54 in86_54 sp86_54 78000.000000
Rwpos86_55 in86_55 sp86_55 78000.000000
Rwpos86_56 in86_56 sp86_56 202000.000000
Rwpos86_57 in86_57 sp86_57 202000.000000
Rwpos86_58 in86_58 sp86_58 78000.000000
Rwpos86_59 in86_59 sp86_59 202000.000000
Rwpos86_60 in86_60 sp86_60 78000.000000
Rwpos86_61 in86_61 sp86_61 202000.000000
Rwpos86_62 in86_62 sp86_62 202000.000000
Rwpos86_63 in86_63 sp86_63 78000.000000
Rwpos86_64 in86_64 sp86_64 202000.000000
Rwpos86_65 in86_65 sp86_65 202000.000000
Rwpos86_66 in86_66 sp86_66 78000.000000
Rwpos86_67 in86_67 sp86_67 78000.000000
Rwpos86_68 in86_68 sp86_68 78000.000000
Rwpos86_69 in86_69 sp86_69 202000.000000
Rwpos86_70 in86_70 sp86_70 78000.000000
Rwpos86_71 in86_71 sp86_71 202000.000000
Rwpos86_72 in86_72 sp86_72 202000.000000
Rwpos86_73 in86_73 sp86_73 78000.000000
Rwpos86_74 in86_74 sp86_74 78000.000000
Rwpos86_75 in86_75 sp86_75 202000.000000
Rwpos86_76 in86_76 sp86_76 78000.000000
Rwpos86_77 in86_77 sp86_77 202000.000000
Rwpos86_78 in86_78 sp86_78 78000.000000
Rwpos86_79 in86_79 sp86_79 78000.000000
Rwpos86_80 in86_80 sp86_80 202000.000000
Rwpos86_81 in86_81 sp86_81 202000.000000
Rwpos86_82 in86_82 sp86_82 202000.000000
Rwpos86_83 in86_83 sp86_83 202000.000000
Rwpos86_84 in86_84 sp86_84 202000.000000
Rwpos87_1 in87_1 sp87_1 202000.000000
Rwpos87_2 in87_2 sp87_2 202000.000000
Rwpos87_3 in87_3 sp87_3 202000.000000
Rwpos87_4 in87_4 sp87_4 78000.000000
Rwpos87_5 in87_5 sp87_5 78000.000000
Rwpos87_6 in87_6 sp87_6 202000.000000
Rwpos87_7 in87_7 sp87_7 78000.000000
Rwpos87_8 in87_8 sp87_8 202000.000000
Rwpos87_9 in87_9 sp87_9 78000.000000
Rwpos87_10 in87_10 sp87_10 202000.000000
Rwpos87_11 in87_11 sp87_11 78000.000000
Rwpos87_12 in87_12 sp87_12 202000.000000
Rwpos87_13 in87_13 sp87_13 78000.000000
Rwpos87_14 in87_14 sp87_14 78000.000000
Rwpos87_15 in87_15 sp87_15 78000.000000
Rwpos87_16 in87_16 sp87_16 78000.000000
Rwpos87_17 in87_17 sp87_17 202000.000000
Rwpos87_18 in87_18 sp87_18 202000.000000
Rwpos87_19 in87_19 sp87_19 202000.000000
Rwpos87_20 in87_20 sp87_20 202000.000000
Rwpos87_21 in87_21 sp87_21 78000.000000
Rwpos87_22 in87_22 sp87_22 202000.000000
Rwpos87_23 in87_23 sp87_23 202000.000000
Rwpos87_24 in87_24 sp87_24 78000.000000
Rwpos87_25 in87_25 sp87_25 78000.000000
Rwpos87_26 in87_26 sp87_26 202000.000000
Rwpos87_27 in87_27 sp87_27 78000.000000
Rwpos87_28 in87_28 sp87_28 78000.000000
Rwpos87_29 in87_29 sp87_29 202000.000000
Rwpos87_30 in87_30 sp87_30 202000.000000
Rwpos87_31 in87_31 sp87_31 202000.000000
Rwpos87_32 in87_32 sp87_32 202000.000000
Rwpos87_33 in87_33 sp87_33 78000.000000
Rwpos87_34 in87_34 sp87_34 202000.000000
Rwpos87_35 in87_35 sp87_35 78000.000000
Rwpos87_36 in87_36 sp87_36 78000.000000
Rwpos87_37 in87_37 sp87_37 78000.000000
Rwpos87_38 in87_38 sp87_38 202000.000000
Rwpos87_39 in87_39 sp87_39 202000.000000
Rwpos87_40 in87_40 sp87_40 202000.000000
Rwpos87_41 in87_41 sp87_41 78000.000000
Rwpos87_42 in87_42 sp87_42 202000.000000
Rwpos87_43 in87_43 sp87_43 202000.000000
Rwpos87_44 in87_44 sp87_44 202000.000000
Rwpos87_45 in87_45 sp87_45 202000.000000
Rwpos87_46 in87_46 sp87_46 78000.000000
Rwpos87_47 in87_47 sp87_47 78000.000000
Rwpos87_48 in87_48 sp87_48 78000.000000
Rwpos87_49 in87_49 sp87_49 78000.000000
Rwpos87_50 in87_50 sp87_50 78000.000000
Rwpos87_51 in87_51 sp87_51 78000.000000
Rwpos87_52 in87_52 sp87_52 78000.000000
Rwpos87_53 in87_53 sp87_53 202000.000000
Rwpos87_54 in87_54 sp87_54 78000.000000
Rwpos87_55 in87_55 sp87_55 202000.000000
Rwpos87_56 in87_56 sp87_56 202000.000000
Rwpos87_57 in87_57 sp87_57 78000.000000
Rwpos87_58 in87_58 sp87_58 202000.000000
Rwpos87_59 in87_59 sp87_59 78000.000000
Rwpos87_60 in87_60 sp87_60 202000.000000
Rwpos87_61 in87_61 sp87_61 202000.000000
Rwpos87_62 in87_62 sp87_62 78000.000000
Rwpos87_63 in87_63 sp87_63 202000.000000
Rwpos87_64 in87_64 sp87_64 202000.000000
Rwpos87_65 in87_65 sp87_65 78000.000000
Rwpos87_66 in87_66 sp87_66 78000.000000
Rwpos87_67 in87_67 sp87_67 78000.000000
Rwpos87_68 in87_68 sp87_68 202000.000000
Rwpos87_69 in87_69 sp87_69 202000.000000
Rwpos87_70 in87_70 sp87_70 78000.000000
Rwpos87_71 in87_71 sp87_71 202000.000000
Rwpos87_72 in87_72 sp87_72 202000.000000
Rwpos87_73 in87_73 sp87_73 202000.000000
Rwpos87_74 in87_74 sp87_74 202000.000000
Rwpos87_75 in87_75 sp87_75 78000.000000
Rwpos87_76 in87_76 sp87_76 78000.000000
Rwpos87_77 in87_77 sp87_77 202000.000000
Rwpos87_78 in87_78 sp87_78 78000.000000
Rwpos87_79 in87_79 sp87_79 202000.000000
Rwpos87_80 in87_80 sp87_80 78000.000000
Rwpos87_81 in87_81 sp87_81 202000.000000
Rwpos87_82 in87_82 sp87_82 78000.000000
Rwpos87_83 in87_83 sp87_83 202000.000000
Rwpos87_84 in87_84 sp87_84 202000.000000
Rwpos88_1 in88_1 sp88_1 202000.000000
Rwpos88_2 in88_2 sp88_2 78000.000000
Rwpos88_3 in88_3 sp88_3 78000.000000
Rwpos88_4 in88_4 sp88_4 202000.000000
Rwpos88_5 in88_5 sp88_5 78000.000000
Rwpos88_6 in88_6 sp88_6 78000.000000
Rwpos88_7 in88_7 sp88_7 78000.000000
Rwpos88_8 in88_8 sp88_8 202000.000000
Rwpos88_9 in88_9 sp88_9 202000.000000
Rwpos88_10 in88_10 sp88_10 202000.000000
Rwpos88_11 in88_11 sp88_11 78000.000000
Rwpos88_12 in88_12 sp88_12 202000.000000
Rwpos88_13 in88_13 sp88_13 202000.000000
Rwpos88_14 in88_14 sp88_14 78000.000000
Rwpos88_15 in88_15 sp88_15 78000.000000
Rwpos88_16 in88_16 sp88_16 78000.000000
Rwpos88_17 in88_17 sp88_17 78000.000000
Rwpos88_18 in88_18 sp88_18 202000.000000
Rwpos88_19 in88_19 sp88_19 78000.000000
Rwpos88_20 in88_20 sp88_20 202000.000000
Rwpos88_21 in88_21 sp88_21 202000.000000
Rwpos88_22 in88_22 sp88_22 78000.000000
Rwpos88_23 in88_23 sp88_23 78000.000000
Rwpos88_24 in88_24 sp88_24 78000.000000
Rwpos88_25 in88_25 sp88_25 78000.000000
Rwpos88_26 in88_26 sp88_26 202000.000000
Rwpos88_27 in88_27 sp88_27 78000.000000
Rwpos88_28 in88_28 sp88_28 202000.000000
Rwpos88_29 in88_29 sp88_29 202000.000000
Rwpos88_30 in88_30 sp88_30 202000.000000
Rwpos88_31 in88_31 sp88_31 202000.000000
Rwpos88_32 in88_32 sp88_32 78000.000000
Rwpos88_33 in88_33 sp88_33 78000.000000
Rwpos88_34 in88_34 sp88_34 202000.000000
Rwpos88_35 in88_35 sp88_35 202000.000000
Rwpos88_36 in88_36 sp88_36 78000.000000
Rwpos88_37 in88_37 sp88_37 202000.000000
Rwpos88_38 in88_38 sp88_38 78000.000000
Rwpos88_39 in88_39 sp88_39 202000.000000
Rwpos88_40 in88_40 sp88_40 78000.000000
Rwpos88_41 in88_41 sp88_41 202000.000000
Rwpos88_42 in88_42 sp88_42 78000.000000
Rwpos88_43 in88_43 sp88_43 202000.000000
Rwpos88_44 in88_44 sp88_44 78000.000000
Rwpos88_45 in88_45 sp88_45 202000.000000
Rwpos88_46 in88_46 sp88_46 78000.000000
Rwpos88_47 in88_47 sp88_47 78000.000000
Rwpos88_48 in88_48 sp88_48 202000.000000
Rwpos88_49 in88_49 sp88_49 202000.000000
Rwpos88_50 in88_50 sp88_50 202000.000000
Rwpos88_51 in88_51 sp88_51 202000.000000
Rwpos88_52 in88_52 sp88_52 202000.000000
Rwpos88_53 in88_53 sp88_53 78000.000000
Rwpos88_54 in88_54 sp88_54 202000.000000
Rwpos88_55 in88_55 sp88_55 78000.000000
Rwpos88_56 in88_56 sp88_56 202000.000000
Rwpos88_57 in88_57 sp88_57 202000.000000
Rwpos88_58 in88_58 sp88_58 78000.000000
Rwpos88_59 in88_59 sp88_59 202000.000000
Rwpos88_60 in88_60 sp88_60 78000.000000
Rwpos88_61 in88_61 sp88_61 202000.000000
Rwpos88_62 in88_62 sp88_62 78000.000000
Rwpos88_63 in88_63 sp88_63 202000.000000
Rwpos88_64 in88_64 sp88_64 202000.000000
Rwpos88_65 in88_65 sp88_65 202000.000000
Rwpos88_66 in88_66 sp88_66 202000.000000
Rwpos88_67 in88_67 sp88_67 78000.000000
Rwpos88_68 in88_68 sp88_68 78000.000000
Rwpos88_69 in88_69 sp88_69 202000.000000
Rwpos88_70 in88_70 sp88_70 202000.000000
Rwpos88_71 in88_71 sp88_71 202000.000000
Rwpos88_72 in88_72 sp88_72 78000.000000
Rwpos88_73 in88_73 sp88_73 202000.000000
Rwpos88_74 in88_74 sp88_74 78000.000000
Rwpos88_75 in88_75 sp88_75 202000.000000
Rwpos88_76 in88_76 sp88_76 202000.000000
Rwpos88_77 in88_77 sp88_77 202000.000000
Rwpos88_78 in88_78 sp88_78 78000.000000
Rwpos88_79 in88_79 sp88_79 202000.000000
Rwpos88_80 in88_80 sp88_80 202000.000000
Rwpos88_81 in88_81 sp88_81 78000.000000
Rwpos88_82 in88_82 sp88_82 202000.000000
Rwpos88_83 in88_83 sp88_83 78000.000000
Rwpos88_84 in88_84 sp88_84 202000.000000
Rwpos89_1 in89_1 sp89_1 202000.000000
Rwpos89_2 in89_2 sp89_2 202000.000000
Rwpos89_3 in89_3 sp89_3 202000.000000
Rwpos89_4 in89_4 sp89_4 202000.000000
Rwpos89_5 in89_5 sp89_5 78000.000000
Rwpos89_6 in89_6 sp89_6 202000.000000
Rwpos89_7 in89_7 sp89_7 78000.000000
Rwpos89_8 in89_8 sp89_8 202000.000000
Rwpos89_9 in89_9 sp89_9 202000.000000
Rwpos89_10 in89_10 sp89_10 78000.000000
Rwpos89_11 in89_11 sp89_11 202000.000000
Rwpos89_12 in89_12 sp89_12 202000.000000
Rwpos89_13 in89_13 sp89_13 78000.000000
Rwpos89_14 in89_14 sp89_14 78000.000000
Rwpos89_15 in89_15 sp89_15 78000.000000
Rwpos89_16 in89_16 sp89_16 202000.000000
Rwpos89_17 in89_17 sp89_17 78000.000000
Rwpos89_18 in89_18 sp89_18 202000.000000
Rwpos89_19 in89_19 sp89_19 202000.000000
Rwpos89_20 in89_20 sp89_20 202000.000000
Rwpos89_21 in89_21 sp89_21 202000.000000
Rwpos89_22 in89_22 sp89_22 78000.000000
Rwpos89_23 in89_23 sp89_23 78000.000000
Rwpos89_24 in89_24 sp89_24 78000.000000
Rwpos89_25 in89_25 sp89_25 78000.000000
Rwpos89_26 in89_26 sp89_26 202000.000000
Rwpos89_27 in89_27 sp89_27 78000.000000
Rwpos89_28 in89_28 sp89_28 202000.000000
Rwpos89_29 in89_29 sp89_29 78000.000000
Rwpos89_30 in89_30 sp89_30 78000.000000
Rwpos89_31 in89_31 sp89_31 78000.000000
Rwpos89_32 in89_32 sp89_32 202000.000000
Rwpos89_33 in89_33 sp89_33 78000.000000
Rwpos89_34 in89_34 sp89_34 202000.000000
Rwpos89_35 in89_35 sp89_35 78000.000000
Rwpos89_36 in89_36 sp89_36 202000.000000
Rwpos89_37 in89_37 sp89_37 202000.000000
Rwpos89_38 in89_38 sp89_38 202000.000000
Rwpos89_39 in89_39 sp89_39 202000.000000
Rwpos89_40 in89_40 sp89_40 78000.000000
Rwpos89_41 in89_41 sp89_41 202000.000000
Rwpos89_42 in89_42 sp89_42 202000.000000
Rwpos89_43 in89_43 sp89_43 78000.000000
Rwpos89_44 in89_44 sp89_44 202000.000000
Rwpos89_45 in89_45 sp89_45 202000.000000
Rwpos89_46 in89_46 sp89_46 78000.000000
Rwpos89_47 in89_47 sp89_47 202000.000000
Rwpos89_48 in89_48 sp89_48 202000.000000
Rwpos89_49 in89_49 sp89_49 202000.000000
Rwpos89_50 in89_50 sp89_50 202000.000000
Rwpos89_51 in89_51 sp89_51 78000.000000
Rwpos89_52 in89_52 sp89_52 202000.000000
Rwpos89_53 in89_53 sp89_53 78000.000000
Rwpos89_54 in89_54 sp89_54 78000.000000
Rwpos89_55 in89_55 sp89_55 202000.000000
Rwpos89_56 in89_56 sp89_56 202000.000000
Rwpos89_57 in89_57 sp89_57 78000.000000
Rwpos89_58 in89_58 sp89_58 78000.000000
Rwpos89_59 in89_59 sp89_59 78000.000000
Rwpos89_60 in89_60 sp89_60 78000.000000
Rwpos89_61 in89_61 sp89_61 202000.000000
Rwpos89_62 in89_62 sp89_62 78000.000000
Rwpos89_63 in89_63 sp89_63 202000.000000
Rwpos89_64 in89_64 sp89_64 202000.000000
Rwpos89_65 in89_65 sp89_65 202000.000000
Rwpos89_66 in89_66 sp89_66 78000.000000
Rwpos89_67 in89_67 sp89_67 78000.000000
Rwpos89_68 in89_68 sp89_68 78000.000000
Rwpos89_69 in89_69 sp89_69 202000.000000
Rwpos89_70 in89_70 sp89_70 78000.000000
Rwpos89_71 in89_71 sp89_71 202000.000000
Rwpos89_72 in89_72 sp89_72 78000.000000
Rwpos89_73 in89_73 sp89_73 78000.000000
Rwpos89_74 in89_74 sp89_74 78000.000000
Rwpos89_75 in89_75 sp89_75 202000.000000
Rwpos89_76 in89_76 sp89_76 202000.000000
Rwpos89_77 in89_77 sp89_77 202000.000000
Rwpos89_78 in89_78 sp89_78 202000.000000
Rwpos89_79 in89_79 sp89_79 202000.000000
Rwpos89_80 in89_80 sp89_80 78000.000000
Rwpos89_81 in89_81 sp89_81 78000.000000
Rwpos89_82 in89_82 sp89_82 202000.000000
Rwpos89_83 in89_83 sp89_83 78000.000000
Rwpos89_84 in89_84 sp89_84 202000.000000
Rwpos90_1 in90_1 sp90_1 202000.000000
Rwpos90_2 in90_2 sp90_2 78000.000000
Rwpos90_3 in90_3 sp90_3 78000.000000
Rwpos90_4 in90_4 sp90_4 78000.000000
Rwpos90_5 in90_5 sp90_5 202000.000000
Rwpos90_6 in90_6 sp90_6 78000.000000
Rwpos90_7 in90_7 sp90_7 202000.000000
Rwpos90_8 in90_8 sp90_8 78000.000000
Rwpos90_9 in90_9 sp90_9 202000.000000
Rwpos90_10 in90_10 sp90_10 78000.000000
Rwpos90_11 in90_11 sp90_11 202000.000000
Rwpos90_12 in90_12 sp90_12 78000.000000
Rwpos90_13 in90_13 sp90_13 78000.000000
Rwpos90_14 in90_14 sp90_14 78000.000000
Rwpos90_15 in90_15 sp90_15 78000.000000
Rwpos90_16 in90_16 sp90_16 202000.000000
Rwpos90_17 in90_17 sp90_17 78000.000000
Rwpos90_18 in90_18 sp90_18 202000.000000
Rwpos90_19 in90_19 sp90_19 202000.000000
Rwpos90_20 in90_20 sp90_20 202000.000000
Rwpos90_21 in90_21 sp90_21 78000.000000
Rwpos90_22 in90_22 sp90_22 78000.000000
Rwpos90_23 in90_23 sp90_23 78000.000000
Rwpos90_24 in90_24 sp90_24 78000.000000
Rwpos90_25 in90_25 sp90_25 78000.000000
Rwpos90_26 in90_26 sp90_26 78000.000000
Rwpos90_27 in90_27 sp90_27 78000.000000
Rwpos90_28 in90_28 sp90_28 202000.000000
Rwpos90_29 in90_29 sp90_29 202000.000000
Rwpos90_30 in90_30 sp90_30 202000.000000
Rwpos90_31 in90_31 sp90_31 78000.000000
Rwpos90_32 in90_32 sp90_32 202000.000000
Rwpos90_33 in90_33 sp90_33 202000.000000
Rwpos90_34 in90_34 sp90_34 202000.000000
Rwpos90_35 in90_35 sp90_35 78000.000000
Rwpos90_36 in90_36 sp90_36 78000.000000
Rwpos90_37 in90_37 sp90_37 202000.000000
Rwpos90_38 in90_38 sp90_38 202000.000000
Rwpos90_39 in90_39 sp90_39 202000.000000
Rwpos90_40 in90_40 sp90_40 202000.000000
Rwpos90_41 in90_41 sp90_41 78000.000000
Rwpos90_42 in90_42 sp90_42 202000.000000
Rwpos90_43 in90_43 sp90_43 78000.000000
Rwpos90_44 in90_44 sp90_44 78000.000000
Rwpos90_45 in90_45 sp90_45 202000.000000
Rwpos90_46 in90_46 sp90_46 78000.000000
Rwpos90_47 in90_47 sp90_47 78000.000000
Rwpos90_48 in90_48 sp90_48 202000.000000
Rwpos90_49 in90_49 sp90_49 202000.000000
Rwpos90_50 in90_50 sp90_50 202000.000000
Rwpos90_51 in90_51 sp90_51 78000.000000
Rwpos90_52 in90_52 sp90_52 202000.000000
Rwpos90_53 in90_53 sp90_53 202000.000000
Rwpos90_54 in90_54 sp90_54 78000.000000
Rwpos90_55 in90_55 sp90_55 202000.000000
Rwpos90_56 in90_56 sp90_56 202000.000000
Rwpos90_57 in90_57 sp90_57 202000.000000
Rwpos90_58 in90_58 sp90_58 78000.000000
Rwpos90_59 in90_59 sp90_59 78000.000000
Rwpos90_60 in90_60 sp90_60 78000.000000
Rwpos90_61 in90_61 sp90_61 78000.000000
Rwpos90_62 in90_62 sp90_62 78000.000000
Rwpos90_63 in90_63 sp90_63 78000.000000
Rwpos90_64 in90_64 sp90_64 202000.000000
Rwpos90_65 in90_65 sp90_65 78000.000000
Rwpos90_66 in90_66 sp90_66 202000.000000
Rwpos90_67 in90_67 sp90_67 78000.000000
Rwpos90_68 in90_68 sp90_68 78000.000000
Rwpos90_69 in90_69 sp90_69 202000.000000
Rwpos90_70 in90_70 sp90_70 78000.000000
Rwpos90_71 in90_71 sp90_71 202000.000000
Rwpos90_72 in90_72 sp90_72 78000.000000
Rwpos90_73 in90_73 sp90_73 78000.000000
Rwpos90_74 in90_74 sp90_74 78000.000000
Rwpos90_75 in90_75 sp90_75 202000.000000
Rwpos90_76 in90_76 sp90_76 78000.000000
Rwpos90_77 in90_77 sp90_77 78000.000000
Rwpos90_78 in90_78 sp90_78 78000.000000
Rwpos90_79 in90_79 sp90_79 202000.000000
Rwpos90_80 in90_80 sp90_80 78000.000000
Rwpos90_81 in90_81 sp90_81 78000.000000
Rwpos90_82 in90_82 sp90_82 78000.000000
Rwpos90_83 in90_83 sp90_83 78000.000000
Rwpos90_84 in90_84 sp90_84 78000.000000
Rwpos91_1 in91_1 sp91_1 78000.000000
Rwpos91_2 in91_2 sp91_2 78000.000000
Rwpos91_3 in91_3 sp91_3 202000.000000
Rwpos91_4 in91_4 sp91_4 202000.000000
Rwpos91_5 in91_5 sp91_5 202000.000000
Rwpos91_6 in91_6 sp91_6 78000.000000
Rwpos91_7 in91_7 sp91_7 78000.000000
Rwpos91_8 in91_8 sp91_8 78000.000000
Rwpos91_9 in91_9 sp91_9 78000.000000
Rwpos91_10 in91_10 sp91_10 78000.000000
Rwpos91_11 in91_11 sp91_11 78000.000000
Rwpos91_12 in91_12 sp91_12 78000.000000
Rwpos91_13 in91_13 sp91_13 202000.000000
Rwpos91_14 in91_14 sp91_14 202000.000000
Rwpos91_15 in91_15 sp91_15 78000.000000
Rwpos91_16 in91_16 sp91_16 78000.000000
Rwpos91_17 in91_17 sp91_17 78000.000000
Rwpos91_18 in91_18 sp91_18 78000.000000
Rwpos91_19 in91_19 sp91_19 78000.000000
Rwpos91_20 in91_20 sp91_20 202000.000000
Rwpos91_21 in91_21 sp91_21 78000.000000
Rwpos91_22 in91_22 sp91_22 78000.000000
Rwpos91_23 in91_23 sp91_23 202000.000000
Rwpos91_24 in91_24 sp91_24 78000.000000
Rwpos91_25 in91_25 sp91_25 78000.000000
Rwpos91_26 in91_26 sp91_26 202000.000000
Rwpos91_27 in91_27 sp91_27 78000.000000
Rwpos91_28 in91_28 sp91_28 78000.000000
Rwpos91_29 in91_29 sp91_29 202000.000000
Rwpos91_30 in91_30 sp91_30 78000.000000
Rwpos91_31 in91_31 sp91_31 202000.000000
Rwpos91_32 in91_32 sp91_32 78000.000000
Rwpos91_33 in91_33 sp91_33 78000.000000
Rwpos91_34 in91_34 sp91_34 202000.000000
Rwpos91_35 in91_35 sp91_35 202000.000000
Rwpos91_36 in91_36 sp91_36 202000.000000
Rwpos91_37 in91_37 sp91_37 78000.000000
Rwpos91_38 in91_38 sp91_38 202000.000000
Rwpos91_39 in91_39 sp91_39 202000.000000
Rwpos91_40 in91_40 sp91_40 78000.000000
Rwpos91_41 in91_41 sp91_41 78000.000000
Rwpos91_42 in91_42 sp91_42 202000.000000
Rwpos91_43 in91_43 sp91_43 78000.000000
Rwpos91_44 in91_44 sp91_44 78000.000000
Rwpos91_45 in91_45 sp91_45 78000.000000
Rwpos91_46 in91_46 sp91_46 202000.000000
Rwpos91_47 in91_47 sp91_47 202000.000000
Rwpos91_48 in91_48 sp91_48 202000.000000
Rwpos91_49 in91_49 sp91_49 202000.000000
Rwpos91_50 in91_50 sp91_50 202000.000000
Rwpos91_51 in91_51 sp91_51 202000.000000
Rwpos91_52 in91_52 sp91_52 202000.000000
Rwpos91_53 in91_53 sp91_53 202000.000000
Rwpos91_54 in91_54 sp91_54 78000.000000
Rwpos91_55 in91_55 sp91_55 78000.000000
Rwpos91_56 in91_56 sp91_56 78000.000000
Rwpos91_57 in91_57 sp91_57 202000.000000
Rwpos91_58 in91_58 sp91_58 78000.000000
Rwpos91_59 in91_59 sp91_59 202000.000000
Rwpos91_60 in91_60 sp91_60 202000.000000
Rwpos91_61 in91_61 sp91_61 78000.000000
Rwpos91_62 in91_62 sp91_62 78000.000000
Rwpos91_63 in91_63 sp91_63 78000.000000
Rwpos91_64 in91_64 sp91_64 202000.000000
Rwpos91_65 in91_65 sp91_65 78000.000000
Rwpos91_66 in91_66 sp91_66 78000.000000
Rwpos91_67 in91_67 sp91_67 202000.000000
Rwpos91_68 in91_68 sp91_68 78000.000000
Rwpos91_69 in91_69 sp91_69 78000.000000
Rwpos91_70 in91_70 sp91_70 202000.000000
Rwpos91_71 in91_71 sp91_71 78000.000000
Rwpos91_72 in91_72 sp91_72 78000.000000
Rwpos91_73 in91_73 sp91_73 78000.000000
Rwpos91_74 in91_74 sp91_74 202000.000000
Rwpos91_75 in91_75 sp91_75 202000.000000
Rwpos91_76 in91_76 sp91_76 202000.000000
Rwpos91_77 in91_77 sp91_77 78000.000000
Rwpos91_78 in91_78 sp91_78 202000.000000
Rwpos91_79 in91_79 sp91_79 202000.000000
Rwpos91_80 in91_80 sp91_80 78000.000000
Rwpos91_81 in91_81 sp91_81 202000.000000
Rwpos91_82 in91_82 sp91_82 78000.000000
Rwpos91_83 in91_83 sp91_83 202000.000000
Rwpos91_84 in91_84 sp91_84 202000.000000
Rwpos92_1 in92_1 sp92_1 202000.000000
Rwpos92_2 in92_2 sp92_2 78000.000000
Rwpos92_3 in92_3 sp92_3 78000.000000
Rwpos92_4 in92_4 sp92_4 202000.000000
Rwpos92_5 in92_5 sp92_5 202000.000000
Rwpos92_6 in92_6 sp92_6 78000.000000
Rwpos92_7 in92_7 sp92_7 78000.000000
Rwpos92_8 in92_8 sp92_8 78000.000000
Rwpos92_9 in92_9 sp92_9 202000.000000
Rwpos92_10 in92_10 sp92_10 202000.000000
Rwpos92_11 in92_11 sp92_11 202000.000000
Rwpos92_12 in92_12 sp92_12 202000.000000
Rwpos92_13 in92_13 sp92_13 202000.000000
Rwpos92_14 in92_14 sp92_14 78000.000000
Rwpos92_15 in92_15 sp92_15 78000.000000
Rwpos92_16 in92_16 sp92_16 202000.000000
Rwpos92_17 in92_17 sp92_17 78000.000000
Rwpos92_18 in92_18 sp92_18 78000.000000
Rwpos92_19 in92_19 sp92_19 202000.000000
Rwpos92_20 in92_20 sp92_20 78000.000000
Rwpos92_21 in92_21 sp92_21 202000.000000
Rwpos92_22 in92_22 sp92_22 202000.000000
Rwpos92_23 in92_23 sp92_23 78000.000000
Rwpos92_24 in92_24 sp92_24 78000.000000
Rwpos92_25 in92_25 sp92_25 78000.000000
Rwpos92_26 in92_26 sp92_26 202000.000000
Rwpos92_27 in92_27 sp92_27 202000.000000
Rwpos92_28 in92_28 sp92_28 78000.000000
Rwpos92_29 in92_29 sp92_29 202000.000000
Rwpos92_30 in92_30 sp92_30 78000.000000
Rwpos92_31 in92_31 sp92_31 202000.000000
Rwpos92_32 in92_32 sp92_32 78000.000000
Rwpos92_33 in92_33 sp92_33 78000.000000
Rwpos92_34 in92_34 sp92_34 202000.000000
Rwpos92_35 in92_35 sp92_35 78000.000000
Rwpos92_36 in92_36 sp92_36 78000.000000
Rwpos92_37 in92_37 sp92_37 202000.000000
Rwpos92_38 in92_38 sp92_38 202000.000000
Rwpos92_39 in92_39 sp92_39 202000.000000
Rwpos92_40 in92_40 sp92_40 202000.000000
Rwpos92_41 in92_41 sp92_41 78000.000000
Rwpos92_42 in92_42 sp92_42 78000.000000
Rwpos92_43 in92_43 sp92_43 202000.000000
Rwpos92_44 in92_44 sp92_44 78000.000000
Rwpos92_45 in92_45 sp92_45 78000.000000
Rwpos92_46 in92_46 sp92_46 78000.000000
Rwpos92_47 in92_47 sp92_47 78000.000000
Rwpos92_48 in92_48 sp92_48 78000.000000
Rwpos92_49 in92_49 sp92_49 202000.000000
Rwpos92_50 in92_50 sp92_50 202000.000000
Rwpos92_51 in92_51 sp92_51 202000.000000
Rwpos92_52 in92_52 sp92_52 202000.000000
Rwpos92_53 in92_53 sp92_53 202000.000000
Rwpos92_54 in92_54 sp92_54 202000.000000
Rwpos92_55 in92_55 sp92_55 78000.000000
Rwpos92_56 in92_56 sp92_56 78000.000000
Rwpos92_57 in92_57 sp92_57 78000.000000
Rwpos92_58 in92_58 sp92_58 78000.000000
Rwpos92_59 in92_59 sp92_59 202000.000000
Rwpos92_60 in92_60 sp92_60 202000.000000
Rwpos92_61 in92_61 sp92_61 78000.000000
Rwpos92_62 in92_62 sp92_62 202000.000000
Rwpos92_63 in92_63 sp92_63 78000.000000
Rwpos92_64 in92_64 sp92_64 202000.000000
Rwpos92_65 in92_65 sp92_65 202000.000000
Rwpos92_66 in92_66 sp92_66 202000.000000
Rwpos92_67 in92_67 sp92_67 202000.000000
Rwpos92_68 in92_68 sp92_68 78000.000000
Rwpos92_69 in92_69 sp92_69 202000.000000
Rwpos92_70 in92_70 sp92_70 78000.000000
Rwpos92_71 in92_71 sp92_71 78000.000000
Rwpos92_72 in92_72 sp92_72 78000.000000
Rwpos92_73 in92_73 sp92_73 202000.000000
Rwpos92_74 in92_74 sp92_74 78000.000000
Rwpos92_75 in92_75 sp92_75 78000.000000
Rwpos92_76 in92_76 sp92_76 78000.000000
Rwpos92_77 in92_77 sp92_77 78000.000000
Rwpos92_78 in92_78 sp92_78 78000.000000
Rwpos92_79 in92_79 sp92_79 78000.000000
Rwpos92_80 in92_80 sp92_80 78000.000000
Rwpos92_81 in92_81 sp92_81 78000.000000
Rwpos92_82 in92_82 sp92_82 78000.000000
Rwpos92_83 in92_83 sp92_83 78000.000000
Rwpos92_84 in92_84 sp92_84 78000.000000
Rwpos93_1 in93_1 sp93_1 78000.000000
Rwpos93_2 in93_2 sp93_2 202000.000000
Rwpos93_3 in93_3 sp93_3 202000.000000
Rwpos93_4 in93_4 sp93_4 202000.000000
Rwpos93_5 in93_5 sp93_5 202000.000000
Rwpos93_6 in93_6 sp93_6 202000.000000
Rwpos93_7 in93_7 sp93_7 78000.000000
Rwpos93_8 in93_8 sp93_8 78000.000000
Rwpos93_9 in93_9 sp93_9 78000.000000
Rwpos93_10 in93_10 sp93_10 78000.000000
Rwpos93_11 in93_11 sp93_11 78000.000000
Rwpos93_12 in93_12 sp93_12 78000.000000
Rwpos93_13 in93_13 sp93_13 78000.000000
Rwpos93_14 in93_14 sp93_14 78000.000000
Rwpos93_15 in93_15 sp93_15 78000.000000
Rwpos93_16 in93_16 sp93_16 78000.000000
Rwpos93_17 in93_17 sp93_17 78000.000000
Rwpos93_18 in93_18 sp93_18 78000.000000
Rwpos93_19 in93_19 sp93_19 202000.000000
Rwpos93_20 in93_20 sp93_20 202000.000000
Rwpos93_21 in93_21 sp93_21 78000.000000
Rwpos93_22 in93_22 sp93_22 202000.000000
Rwpos93_23 in93_23 sp93_23 202000.000000
Rwpos93_24 in93_24 sp93_24 78000.000000
Rwpos93_25 in93_25 sp93_25 202000.000000
Rwpos93_26 in93_26 sp93_26 78000.000000
Rwpos93_27 in93_27 sp93_27 78000.000000
Rwpos93_28 in93_28 sp93_28 78000.000000
Rwpos93_29 in93_29 sp93_29 202000.000000
Rwpos93_30 in93_30 sp93_30 202000.000000
Rwpos93_31 in93_31 sp93_31 78000.000000
Rwpos93_32 in93_32 sp93_32 78000.000000
Rwpos93_33 in93_33 sp93_33 202000.000000
Rwpos93_34 in93_34 sp93_34 78000.000000
Rwpos93_35 in93_35 sp93_35 202000.000000
Rwpos93_36 in93_36 sp93_36 78000.000000
Rwpos93_37 in93_37 sp93_37 78000.000000
Rwpos93_38 in93_38 sp93_38 202000.000000
Rwpos93_39 in93_39 sp93_39 78000.000000
Rwpos93_40 in93_40 sp93_40 202000.000000
Rwpos93_41 in93_41 sp93_41 202000.000000
Rwpos93_42 in93_42 sp93_42 202000.000000
Rwpos93_43 in93_43 sp93_43 78000.000000
Rwpos93_44 in93_44 sp93_44 78000.000000
Rwpos93_45 in93_45 sp93_45 202000.000000
Rwpos93_46 in93_46 sp93_46 78000.000000
Rwpos93_47 in93_47 sp93_47 202000.000000
Rwpos93_48 in93_48 sp93_48 78000.000000
Rwpos93_49 in93_49 sp93_49 202000.000000
Rwpos93_50 in93_50 sp93_50 78000.000000
Rwpos93_51 in93_51 sp93_51 202000.000000
Rwpos93_52 in93_52 sp93_52 78000.000000
Rwpos93_53 in93_53 sp93_53 78000.000000
Rwpos93_54 in93_54 sp93_54 78000.000000
Rwpos93_55 in93_55 sp93_55 78000.000000
Rwpos93_56 in93_56 sp93_56 202000.000000
Rwpos93_57 in93_57 sp93_57 202000.000000
Rwpos93_58 in93_58 sp93_58 202000.000000
Rwpos93_59 in93_59 sp93_59 78000.000000
Rwpos93_60 in93_60 sp93_60 78000.000000
Rwpos93_61 in93_61 sp93_61 78000.000000
Rwpos93_62 in93_62 sp93_62 78000.000000
Rwpos93_63 in93_63 sp93_63 78000.000000
Rwpos93_64 in93_64 sp93_64 78000.000000
Rwpos93_65 in93_65 sp93_65 202000.000000
Rwpos93_66 in93_66 sp93_66 78000.000000
Rwpos93_67 in93_67 sp93_67 78000.000000
Rwpos93_68 in93_68 sp93_68 78000.000000
Rwpos93_69 in93_69 sp93_69 78000.000000
Rwpos93_70 in93_70 sp93_70 202000.000000
Rwpos93_71 in93_71 sp93_71 78000.000000
Rwpos93_72 in93_72 sp93_72 78000.000000
Rwpos93_73 in93_73 sp93_73 78000.000000
Rwpos93_74 in93_74 sp93_74 202000.000000
Rwpos93_75 in93_75 sp93_75 202000.000000
Rwpos93_76 in93_76 sp93_76 78000.000000
Rwpos93_77 in93_77 sp93_77 202000.000000
Rwpos93_78 in93_78 sp93_78 202000.000000
Rwpos93_79 in93_79 sp93_79 78000.000000
Rwpos93_80 in93_80 sp93_80 78000.000000
Rwpos93_81 in93_81 sp93_81 202000.000000
Rwpos93_82 in93_82 sp93_82 78000.000000
Rwpos93_83 in93_83 sp93_83 202000.000000
Rwpos93_84 in93_84 sp93_84 202000.000000
Rwpos94_1 in94_1 sp94_1 202000.000000
Rwpos94_2 in94_2 sp94_2 202000.000000
Rwpos94_3 in94_3 sp94_3 78000.000000
Rwpos94_4 in94_4 sp94_4 78000.000000
Rwpos94_5 in94_5 sp94_5 78000.000000
Rwpos94_6 in94_6 sp94_6 78000.000000
Rwpos94_7 in94_7 sp94_7 202000.000000
Rwpos94_8 in94_8 sp94_8 202000.000000
Rwpos94_9 in94_9 sp94_9 78000.000000
Rwpos94_10 in94_10 sp94_10 78000.000000
Rwpos94_11 in94_11 sp94_11 78000.000000
Rwpos94_12 in94_12 sp94_12 78000.000000
Rwpos94_13 in94_13 sp94_13 202000.000000
Rwpos94_14 in94_14 sp94_14 78000.000000
Rwpos94_15 in94_15 sp94_15 78000.000000
Rwpos94_16 in94_16 sp94_16 202000.000000
Rwpos94_17 in94_17 sp94_17 202000.000000
Rwpos94_18 in94_18 sp94_18 78000.000000
Rwpos94_19 in94_19 sp94_19 78000.000000
Rwpos94_20 in94_20 sp94_20 202000.000000
Rwpos94_21 in94_21 sp94_21 78000.000000
Rwpos94_22 in94_22 sp94_22 202000.000000
Rwpos94_23 in94_23 sp94_23 202000.000000
Rwpos94_24 in94_24 sp94_24 78000.000000
Rwpos94_25 in94_25 sp94_25 202000.000000
Rwpos94_26 in94_26 sp94_26 78000.000000
Rwpos94_27 in94_27 sp94_27 202000.000000
Rwpos94_28 in94_28 sp94_28 202000.000000
Rwpos94_29 in94_29 sp94_29 78000.000000
Rwpos94_30 in94_30 sp94_30 78000.000000
Rwpos94_31 in94_31 sp94_31 78000.000000
Rwpos94_32 in94_32 sp94_32 78000.000000
Rwpos94_33 in94_33 sp94_33 202000.000000
Rwpos94_34 in94_34 sp94_34 78000.000000
Rwpos94_35 in94_35 sp94_35 202000.000000
Rwpos94_36 in94_36 sp94_36 78000.000000
Rwpos94_37 in94_37 sp94_37 78000.000000
Rwpos94_38 in94_38 sp94_38 78000.000000
Rwpos94_39 in94_39 sp94_39 78000.000000
Rwpos94_40 in94_40 sp94_40 202000.000000
Rwpos94_41 in94_41 sp94_41 202000.000000
Rwpos94_42 in94_42 sp94_42 202000.000000
Rwpos94_43 in94_43 sp94_43 78000.000000
Rwpos94_44 in94_44 sp94_44 202000.000000
Rwpos94_45 in94_45 sp94_45 202000.000000
Rwpos94_46 in94_46 sp94_46 78000.000000
Rwpos94_47 in94_47 sp94_47 78000.000000
Rwpos94_48 in94_48 sp94_48 202000.000000
Rwpos94_49 in94_49 sp94_49 202000.000000
Rwpos94_50 in94_50 sp94_50 202000.000000
Rwpos94_51 in94_51 sp94_51 202000.000000
Rwpos94_52 in94_52 sp94_52 78000.000000
Rwpos94_53 in94_53 sp94_53 202000.000000
Rwpos94_54 in94_54 sp94_54 202000.000000
Rwpos94_55 in94_55 sp94_55 78000.000000
Rwpos94_56 in94_56 sp94_56 78000.000000
Rwpos94_57 in94_57 sp94_57 78000.000000
Rwpos94_58 in94_58 sp94_58 202000.000000
Rwpos94_59 in94_59 sp94_59 78000.000000
Rwpos94_60 in94_60 sp94_60 78000.000000
Rwpos94_61 in94_61 sp94_61 78000.000000
Rwpos94_62 in94_62 sp94_62 202000.000000
Rwpos94_63 in94_63 sp94_63 78000.000000
Rwpos94_64 in94_64 sp94_64 78000.000000
Rwpos94_65 in94_65 sp94_65 78000.000000
Rwpos94_66 in94_66 sp94_66 202000.000000
Rwpos94_67 in94_67 sp94_67 78000.000000
Rwpos94_68 in94_68 sp94_68 78000.000000
Rwpos94_69 in94_69 sp94_69 78000.000000
Rwpos94_70 in94_70 sp94_70 78000.000000
Rwpos94_71 in94_71 sp94_71 78000.000000
Rwpos94_72 in94_72 sp94_72 202000.000000
Rwpos94_73 in94_73 sp94_73 78000.000000
Rwpos94_74 in94_74 sp94_74 78000.000000
Rwpos94_75 in94_75 sp94_75 78000.000000
Rwpos94_76 in94_76 sp94_76 78000.000000
Rwpos94_77 in94_77 sp94_77 78000.000000
Rwpos94_78 in94_78 sp94_78 78000.000000
Rwpos94_79 in94_79 sp94_79 78000.000000
Rwpos94_80 in94_80 sp94_80 202000.000000
Rwpos94_81 in94_81 sp94_81 202000.000000
Rwpos94_82 in94_82 sp94_82 78000.000000
Rwpos94_83 in94_83 sp94_83 202000.000000
Rwpos94_84 in94_84 sp94_84 202000.000000
Rwpos95_1 in95_1 sp95_1 202000.000000
Rwpos95_2 in95_2 sp95_2 78000.000000
Rwpos95_3 in95_3 sp95_3 78000.000000
Rwpos95_4 in95_4 sp95_4 78000.000000
Rwpos95_5 in95_5 sp95_5 202000.000000
Rwpos95_6 in95_6 sp95_6 202000.000000
Rwpos95_7 in95_7 sp95_7 78000.000000
Rwpos95_8 in95_8 sp95_8 78000.000000
Rwpos95_9 in95_9 sp95_9 78000.000000
Rwpos95_10 in95_10 sp95_10 202000.000000
Rwpos95_11 in95_11 sp95_11 202000.000000
Rwpos95_12 in95_12 sp95_12 78000.000000
Rwpos95_13 in95_13 sp95_13 78000.000000
Rwpos95_14 in95_14 sp95_14 202000.000000
Rwpos95_15 in95_15 sp95_15 78000.000000
Rwpos95_16 in95_16 sp95_16 78000.000000
Rwpos95_17 in95_17 sp95_17 202000.000000
Rwpos95_18 in95_18 sp95_18 78000.000000
Rwpos95_19 in95_19 sp95_19 202000.000000
Rwpos95_20 in95_20 sp95_20 78000.000000
Rwpos95_21 in95_21 sp95_21 78000.000000
Rwpos95_22 in95_22 sp95_22 78000.000000
Rwpos95_23 in95_23 sp95_23 202000.000000
Rwpos95_24 in95_24 sp95_24 78000.000000
Rwpos95_25 in95_25 sp95_25 202000.000000
Rwpos95_26 in95_26 sp95_26 78000.000000
Rwpos95_27 in95_27 sp95_27 78000.000000
Rwpos95_28 in95_28 sp95_28 78000.000000
Rwpos95_29 in95_29 sp95_29 78000.000000
Rwpos95_30 in95_30 sp95_30 202000.000000
Rwpos95_31 in95_31 sp95_31 202000.000000
Rwpos95_32 in95_32 sp95_32 202000.000000
Rwpos95_33 in95_33 sp95_33 78000.000000
Rwpos95_34 in95_34 sp95_34 78000.000000
Rwpos95_35 in95_35 sp95_35 78000.000000
Rwpos95_36 in95_36 sp95_36 202000.000000
Rwpos95_37 in95_37 sp95_37 78000.000000
Rwpos95_38 in95_38 sp95_38 78000.000000
Rwpos95_39 in95_39 sp95_39 202000.000000
Rwpos95_40 in95_40 sp95_40 202000.000000
Rwpos95_41 in95_41 sp95_41 202000.000000
Rwpos95_42 in95_42 sp95_42 78000.000000
Rwpos95_43 in95_43 sp95_43 202000.000000
Rwpos95_44 in95_44 sp95_44 202000.000000
Rwpos95_45 in95_45 sp95_45 202000.000000
Rwpos95_46 in95_46 sp95_46 78000.000000
Rwpos95_47 in95_47 sp95_47 202000.000000
Rwpos95_48 in95_48 sp95_48 202000.000000
Rwpos95_49 in95_49 sp95_49 78000.000000
Rwpos95_50 in95_50 sp95_50 78000.000000
Rwpos95_51 in95_51 sp95_51 78000.000000
Rwpos95_52 in95_52 sp95_52 78000.000000
Rwpos95_53 in95_53 sp95_53 78000.000000
Rwpos95_54 in95_54 sp95_54 202000.000000
Rwpos95_55 in95_55 sp95_55 202000.000000
Rwpos95_56 in95_56 sp95_56 78000.000000
Rwpos95_57 in95_57 sp95_57 78000.000000
Rwpos95_58 in95_58 sp95_58 202000.000000
Rwpos95_59 in95_59 sp95_59 78000.000000
Rwpos95_60 in95_60 sp95_60 78000.000000
Rwpos95_61 in95_61 sp95_61 78000.000000
Rwpos95_62 in95_62 sp95_62 202000.000000
Rwpos95_63 in95_63 sp95_63 78000.000000
Rwpos95_64 in95_64 sp95_64 78000.000000
Rwpos95_65 in95_65 sp95_65 78000.000000
Rwpos95_66 in95_66 sp95_66 78000.000000
Rwpos95_67 in95_67 sp95_67 202000.000000
Rwpos95_68 in95_68 sp95_68 202000.000000
Rwpos95_69 in95_69 sp95_69 78000.000000
Rwpos95_70 in95_70 sp95_70 78000.000000
Rwpos95_71 in95_71 sp95_71 78000.000000
Rwpos95_72 in95_72 sp95_72 78000.000000
Rwpos95_73 in95_73 sp95_73 202000.000000
Rwpos95_74 in95_74 sp95_74 78000.000000
Rwpos95_75 in95_75 sp95_75 78000.000000
Rwpos95_76 in95_76 sp95_76 202000.000000
Rwpos95_77 in95_77 sp95_77 202000.000000
Rwpos95_78 in95_78 sp95_78 78000.000000
Rwpos95_79 in95_79 sp95_79 202000.000000
Rwpos95_80 in95_80 sp95_80 78000.000000
Rwpos95_81 in95_81 sp95_81 202000.000000
Rwpos95_82 in95_82 sp95_82 78000.000000
Rwpos95_83 in95_83 sp95_83 202000.000000
Rwpos95_84 in95_84 sp95_84 202000.000000
Rwpos96_1 in96_1 sp96_1 78000.000000
Rwpos96_2 in96_2 sp96_2 78000.000000
Rwpos96_3 in96_3 sp96_3 78000.000000
Rwpos96_4 in96_4 sp96_4 202000.000000
Rwpos96_5 in96_5 sp96_5 78000.000000
Rwpos96_6 in96_6 sp96_6 78000.000000
Rwpos96_7 in96_7 sp96_7 78000.000000
Rwpos96_8 in96_8 sp96_8 202000.000000
Rwpos96_9 in96_9 sp96_9 202000.000000
Rwpos96_10 in96_10 sp96_10 202000.000000
Rwpos96_11 in96_11 sp96_11 202000.000000
Rwpos96_12 in96_12 sp96_12 202000.000000
Rwpos96_13 in96_13 sp96_13 78000.000000
Rwpos96_14 in96_14 sp96_14 78000.000000
Rwpos96_15 in96_15 sp96_15 78000.000000
Rwpos96_16 in96_16 sp96_16 202000.000000
Rwpos96_17 in96_17 sp96_17 202000.000000
Rwpos96_18 in96_18 sp96_18 202000.000000
Rwpos96_19 in96_19 sp96_19 78000.000000
Rwpos96_20 in96_20 sp96_20 202000.000000
Rwpos96_21 in96_21 sp96_21 78000.000000
Rwpos96_22 in96_22 sp96_22 78000.000000
Rwpos96_23 in96_23 sp96_23 202000.000000
Rwpos96_24 in96_24 sp96_24 78000.000000
Rwpos96_25 in96_25 sp96_25 202000.000000
Rwpos96_26 in96_26 sp96_26 78000.000000
Rwpos96_27 in96_27 sp96_27 78000.000000
Rwpos96_28 in96_28 sp96_28 78000.000000
Rwpos96_29 in96_29 sp96_29 78000.000000
Rwpos96_30 in96_30 sp96_30 202000.000000
Rwpos96_31 in96_31 sp96_31 202000.000000
Rwpos96_32 in96_32 sp96_32 202000.000000
Rwpos96_33 in96_33 sp96_33 78000.000000
Rwpos96_34 in96_34 sp96_34 202000.000000
Rwpos96_35 in96_35 sp96_35 78000.000000
Rwpos96_36 in96_36 sp96_36 202000.000000
Rwpos96_37 in96_37 sp96_37 202000.000000
Rwpos96_38 in96_38 sp96_38 78000.000000
Rwpos96_39 in96_39 sp96_39 78000.000000
Rwpos96_40 in96_40 sp96_40 78000.000000
Rwpos96_41 in96_41 sp96_41 78000.000000
Rwpos96_42 in96_42 sp96_42 78000.000000
Rwpos96_43 in96_43 sp96_43 202000.000000
Rwpos96_44 in96_44 sp96_44 78000.000000
Rwpos96_45 in96_45 sp96_45 202000.000000
Rwpos96_46 in96_46 sp96_46 202000.000000
Rwpos96_47 in96_47 sp96_47 78000.000000
Rwpos96_48 in96_48 sp96_48 78000.000000
Rwpos96_49 in96_49 sp96_49 78000.000000
Rwpos96_50 in96_50 sp96_50 78000.000000
Rwpos96_51 in96_51 sp96_51 78000.000000
Rwpos96_52 in96_52 sp96_52 78000.000000
Rwpos96_53 in96_53 sp96_53 202000.000000
Rwpos96_54 in96_54 sp96_54 78000.000000
Rwpos96_55 in96_55 sp96_55 78000.000000
Rwpos96_56 in96_56 sp96_56 202000.000000
Rwpos96_57 in96_57 sp96_57 78000.000000
Rwpos96_58 in96_58 sp96_58 202000.000000
Rwpos96_59 in96_59 sp96_59 202000.000000
Rwpos96_60 in96_60 sp96_60 78000.000000
Rwpos96_61 in96_61 sp96_61 202000.000000
Rwpos96_62 in96_62 sp96_62 202000.000000
Rwpos96_63 in96_63 sp96_63 202000.000000
Rwpos96_64 in96_64 sp96_64 78000.000000
Rwpos96_65 in96_65 sp96_65 78000.000000
Rwpos96_66 in96_66 sp96_66 202000.000000
Rwpos96_67 in96_67 sp96_67 78000.000000
Rwpos96_68 in96_68 sp96_68 202000.000000
Rwpos96_69 in96_69 sp96_69 202000.000000
Rwpos96_70 in96_70 sp96_70 202000.000000
Rwpos96_71 in96_71 sp96_71 202000.000000
Rwpos96_72 in96_72 sp96_72 78000.000000
Rwpos96_73 in96_73 sp96_73 202000.000000
Rwpos96_74 in96_74 sp96_74 78000.000000
Rwpos96_75 in96_75 sp96_75 78000.000000
Rwpos96_76 in96_76 sp96_76 78000.000000
Rwpos96_77 in96_77 sp96_77 202000.000000
Rwpos96_78 in96_78 sp96_78 78000.000000
Rwpos96_79 in96_79 sp96_79 202000.000000
Rwpos96_80 in96_80 sp96_80 202000.000000
Rwpos96_81 in96_81 sp96_81 78000.000000
Rwpos96_82 in96_82 sp96_82 202000.000000
Rwpos96_83 in96_83 sp96_83 78000.000000
Rwpos96_84 in96_84 sp96_84 78000.000000
Rwpos97_1 in97_1 sp97_1 202000.000000
Rwpos97_2 in97_2 sp97_2 78000.000000
Rwpos97_3 in97_3 sp97_3 202000.000000
Rwpos97_4 in97_4 sp97_4 78000.000000
Rwpos97_5 in97_5 sp97_5 202000.000000
Rwpos97_6 in97_6 sp97_6 78000.000000
Rwpos97_7 in97_7 sp97_7 78000.000000
Rwpos97_8 in97_8 sp97_8 78000.000000
Rwpos97_9 in97_9 sp97_9 78000.000000
Rwpos97_10 in97_10 sp97_10 202000.000000
Rwpos97_11 in97_11 sp97_11 202000.000000
Rwpos97_12 in97_12 sp97_12 78000.000000
Rwpos97_13 in97_13 sp97_13 202000.000000
Rwpos97_14 in97_14 sp97_14 202000.000000
Rwpos97_15 in97_15 sp97_15 78000.000000
Rwpos97_16 in97_16 sp97_16 78000.000000
Rwpos97_17 in97_17 sp97_17 78000.000000
Rwpos97_18 in97_18 sp97_18 202000.000000
Rwpos97_19 in97_19 sp97_19 78000.000000
Rwpos97_20 in97_20 sp97_20 202000.000000
Rwpos97_21 in97_21 sp97_21 78000.000000
Rwpos97_22 in97_22 sp97_22 78000.000000
Rwpos97_23 in97_23 sp97_23 78000.000000
Rwpos97_24 in97_24 sp97_24 202000.000000
Rwpos97_25 in97_25 sp97_25 78000.000000
Rwpos97_26 in97_26 sp97_26 78000.000000
Rwpos97_27 in97_27 sp97_27 78000.000000
Rwpos97_28 in97_28 sp97_28 202000.000000
Rwpos97_29 in97_29 sp97_29 202000.000000
Rwpos97_30 in97_30 sp97_30 78000.000000
Rwpos97_31 in97_31 sp97_31 78000.000000
Rwpos97_32 in97_32 sp97_32 202000.000000
Rwpos97_33 in97_33 sp97_33 202000.000000
Rwpos97_34 in97_34 sp97_34 202000.000000
Rwpos97_35 in97_35 sp97_35 202000.000000
Rwpos97_36 in97_36 sp97_36 202000.000000
Rwpos97_37 in97_37 sp97_37 202000.000000
Rwpos97_38 in97_38 sp97_38 202000.000000
Rwpos97_39 in97_39 sp97_39 202000.000000
Rwpos97_40 in97_40 sp97_40 202000.000000
Rwpos97_41 in97_41 sp97_41 78000.000000
Rwpos97_42 in97_42 sp97_42 202000.000000
Rwpos97_43 in97_43 sp97_43 78000.000000
Rwpos97_44 in97_44 sp97_44 78000.000000
Rwpos97_45 in97_45 sp97_45 78000.000000
Rwpos97_46 in97_46 sp97_46 202000.000000
Rwpos97_47 in97_47 sp97_47 202000.000000
Rwpos97_48 in97_48 sp97_48 202000.000000
Rwpos97_49 in97_49 sp97_49 78000.000000
Rwpos97_50 in97_50 sp97_50 202000.000000
Rwpos97_51 in97_51 sp97_51 202000.000000
Rwpos97_52 in97_52 sp97_52 78000.000000
Rwpos97_53 in97_53 sp97_53 202000.000000
Rwpos97_54 in97_54 sp97_54 78000.000000
Rwpos97_55 in97_55 sp97_55 202000.000000
Rwpos97_56 in97_56 sp97_56 78000.000000
Rwpos97_57 in97_57 sp97_57 202000.000000
Rwpos97_58 in97_58 sp97_58 78000.000000
Rwpos97_59 in97_59 sp97_59 202000.000000
Rwpos97_60 in97_60 sp97_60 78000.000000
Rwpos97_61 in97_61 sp97_61 78000.000000
Rwpos97_62 in97_62 sp97_62 202000.000000
Rwpos97_63 in97_63 sp97_63 78000.000000
Rwpos97_64 in97_64 sp97_64 202000.000000
Rwpos97_65 in97_65 sp97_65 78000.000000
Rwpos97_66 in97_66 sp97_66 78000.000000
Rwpos97_67 in97_67 sp97_67 202000.000000
Rwpos97_68 in97_68 sp97_68 78000.000000
Rwpos97_69 in97_69 sp97_69 78000.000000
Rwpos97_70 in97_70 sp97_70 78000.000000
Rwpos97_71 in97_71 sp97_71 78000.000000
Rwpos97_72 in97_72 sp97_72 78000.000000
Rwpos97_73 in97_73 sp97_73 78000.000000
Rwpos97_74 in97_74 sp97_74 78000.000000
Rwpos97_75 in97_75 sp97_75 202000.000000
Rwpos97_76 in97_76 sp97_76 78000.000000
Rwpos97_77 in97_77 sp97_77 78000.000000
Rwpos97_78 in97_78 sp97_78 78000.000000
Rwpos97_79 in97_79 sp97_79 78000.000000
Rwpos97_80 in97_80 sp97_80 202000.000000
Rwpos97_81 in97_81 sp97_81 78000.000000
Rwpos97_82 in97_82 sp97_82 78000.000000
Rwpos97_83 in97_83 sp97_83 78000.000000
Rwpos97_84 in97_84 sp97_84 78000.000000
Rwpos98_1 in98_1 sp98_1 78000.000000
Rwpos98_2 in98_2 sp98_2 78000.000000
Rwpos98_3 in98_3 sp98_3 78000.000000
Rwpos98_4 in98_4 sp98_4 78000.000000
Rwpos98_5 in98_5 sp98_5 78000.000000
Rwpos98_6 in98_6 sp98_6 202000.000000
Rwpos98_7 in98_7 sp98_7 202000.000000
Rwpos98_8 in98_8 sp98_8 78000.000000
Rwpos98_9 in98_9 sp98_9 78000.000000
Rwpos98_10 in98_10 sp98_10 78000.000000
Rwpos98_11 in98_11 sp98_11 78000.000000
Rwpos98_12 in98_12 sp98_12 78000.000000
Rwpos98_13 in98_13 sp98_13 78000.000000
Rwpos98_14 in98_14 sp98_14 202000.000000
Rwpos98_15 in98_15 sp98_15 202000.000000
Rwpos98_16 in98_16 sp98_16 202000.000000
Rwpos98_17 in98_17 sp98_17 78000.000000
Rwpos98_18 in98_18 sp98_18 78000.000000
Rwpos98_19 in98_19 sp98_19 202000.000000
Rwpos98_20 in98_20 sp98_20 202000.000000
Rwpos98_21 in98_21 sp98_21 202000.000000
Rwpos98_22 in98_22 sp98_22 202000.000000
Rwpos98_23 in98_23 sp98_23 202000.000000
Rwpos98_24 in98_24 sp98_24 78000.000000
Rwpos98_25 in98_25 sp98_25 78000.000000
Rwpos98_26 in98_26 sp98_26 78000.000000
Rwpos98_27 in98_27 sp98_27 78000.000000
Rwpos98_28 in98_28 sp98_28 202000.000000
Rwpos98_29 in98_29 sp98_29 202000.000000
Rwpos98_30 in98_30 sp98_30 78000.000000
Rwpos98_31 in98_31 sp98_31 202000.000000
Rwpos98_32 in98_32 sp98_32 78000.000000
Rwpos98_33 in98_33 sp98_33 202000.000000
Rwpos98_34 in98_34 sp98_34 78000.000000
Rwpos98_35 in98_35 sp98_35 202000.000000
Rwpos98_36 in98_36 sp98_36 78000.000000
Rwpos98_37 in98_37 sp98_37 202000.000000
Rwpos98_38 in98_38 sp98_38 202000.000000
Rwpos98_39 in98_39 sp98_39 202000.000000
Rwpos98_40 in98_40 sp98_40 202000.000000
Rwpos98_41 in98_41 sp98_41 202000.000000
Rwpos98_42 in98_42 sp98_42 202000.000000
Rwpos98_43 in98_43 sp98_43 202000.000000
Rwpos98_44 in98_44 sp98_44 78000.000000
Rwpos98_45 in98_45 sp98_45 202000.000000
Rwpos98_46 in98_46 sp98_46 202000.000000
Rwpos98_47 in98_47 sp98_47 78000.000000
Rwpos98_48 in98_48 sp98_48 78000.000000
Rwpos98_49 in98_49 sp98_49 78000.000000
Rwpos98_50 in98_50 sp98_50 202000.000000
Rwpos98_51 in98_51 sp98_51 202000.000000
Rwpos98_52 in98_52 sp98_52 202000.000000
Rwpos98_53 in98_53 sp98_53 202000.000000
Rwpos98_54 in98_54 sp98_54 202000.000000
Rwpos98_55 in98_55 sp98_55 202000.000000
Rwpos98_56 in98_56 sp98_56 78000.000000
Rwpos98_57 in98_57 sp98_57 78000.000000
Rwpos98_58 in98_58 sp98_58 202000.000000
Rwpos98_59 in98_59 sp98_59 78000.000000
Rwpos98_60 in98_60 sp98_60 78000.000000
Rwpos98_61 in98_61 sp98_61 202000.000000
Rwpos98_62 in98_62 sp98_62 78000.000000
Rwpos98_63 in98_63 sp98_63 78000.000000
Rwpos98_64 in98_64 sp98_64 78000.000000
Rwpos98_65 in98_65 sp98_65 202000.000000
Rwpos98_66 in98_66 sp98_66 78000.000000
Rwpos98_67 in98_67 sp98_67 202000.000000
Rwpos98_68 in98_68 sp98_68 78000.000000
Rwpos98_69 in98_69 sp98_69 78000.000000
Rwpos98_70 in98_70 sp98_70 78000.000000
Rwpos98_71 in98_71 sp98_71 78000.000000
Rwpos98_72 in98_72 sp98_72 78000.000000
Rwpos98_73 in98_73 sp98_73 78000.000000
Rwpos98_74 in98_74 sp98_74 78000.000000
Rwpos98_75 in98_75 sp98_75 202000.000000
Rwpos98_76 in98_76 sp98_76 78000.000000
Rwpos98_77 in98_77 sp98_77 202000.000000
Rwpos98_78 in98_78 sp98_78 78000.000000
Rwpos98_79 in98_79 sp98_79 78000.000000
Rwpos98_80 in98_80 sp98_80 202000.000000
Rwpos98_81 in98_81 sp98_81 78000.000000
Rwpos98_82 in98_82 sp98_82 78000.000000
Rwpos98_83 in98_83 sp98_83 202000.000000
Rwpos98_84 in98_84 sp98_84 202000.000000
Rwpos99_1 in99_1 sp99_1 78000.000000
Rwpos99_2 in99_2 sp99_2 78000.000000
Rwpos99_3 in99_3 sp99_3 202000.000000
Rwpos99_4 in99_4 sp99_4 78000.000000
Rwpos99_5 in99_5 sp99_5 78000.000000
Rwpos99_6 in99_6 sp99_6 78000.000000
Rwpos99_7 in99_7 sp99_7 202000.000000
Rwpos99_8 in99_8 sp99_8 202000.000000
Rwpos99_9 in99_9 sp99_9 78000.000000
Rwpos99_10 in99_10 sp99_10 78000.000000
Rwpos99_11 in99_11 sp99_11 78000.000000
Rwpos99_12 in99_12 sp99_12 78000.000000
Rwpos99_13 in99_13 sp99_13 78000.000000
Rwpos99_14 in99_14 sp99_14 78000.000000
Rwpos99_15 in99_15 sp99_15 202000.000000
Rwpos99_16 in99_16 sp99_16 78000.000000
Rwpos99_17 in99_17 sp99_17 78000.000000
Rwpos99_18 in99_18 sp99_18 78000.000000
Rwpos99_19 in99_19 sp99_19 78000.000000
Rwpos99_20 in99_20 sp99_20 202000.000000
Rwpos99_21 in99_21 sp99_21 78000.000000
Rwpos99_22 in99_22 sp99_22 78000.000000
Rwpos99_23 in99_23 sp99_23 78000.000000
Rwpos99_24 in99_24 sp99_24 202000.000000
Rwpos99_25 in99_25 sp99_25 78000.000000
Rwpos99_26 in99_26 sp99_26 78000.000000
Rwpos99_27 in99_27 sp99_27 78000.000000
Rwpos99_28 in99_28 sp99_28 78000.000000
Rwpos99_29 in99_29 sp99_29 78000.000000
Rwpos99_30 in99_30 sp99_30 202000.000000
Rwpos99_31 in99_31 sp99_31 78000.000000
Rwpos99_32 in99_32 sp99_32 78000.000000
Rwpos99_33 in99_33 sp99_33 202000.000000
Rwpos99_34 in99_34 sp99_34 78000.000000
Rwpos99_35 in99_35 sp99_35 202000.000000
Rwpos99_36 in99_36 sp99_36 202000.000000
Rwpos99_37 in99_37 sp99_37 202000.000000
Rwpos99_38 in99_38 sp99_38 202000.000000
Rwpos99_39 in99_39 sp99_39 78000.000000
Rwpos99_40 in99_40 sp99_40 78000.000000
Rwpos99_41 in99_41 sp99_41 202000.000000
Rwpos99_42 in99_42 sp99_42 202000.000000
Rwpos99_43 in99_43 sp99_43 202000.000000
Rwpos99_44 in99_44 sp99_44 78000.000000
Rwpos99_45 in99_45 sp99_45 78000.000000
Rwpos99_46 in99_46 sp99_46 78000.000000
Rwpos99_47 in99_47 sp99_47 78000.000000
Rwpos99_48 in99_48 sp99_48 202000.000000
Rwpos99_49 in99_49 sp99_49 202000.000000
Rwpos99_50 in99_50 sp99_50 202000.000000
Rwpos99_51 in99_51 sp99_51 78000.000000
Rwpos99_52 in99_52 sp99_52 202000.000000
Rwpos99_53 in99_53 sp99_53 78000.000000
Rwpos99_54 in99_54 sp99_54 78000.000000
Rwpos99_55 in99_55 sp99_55 202000.000000
Rwpos99_56 in99_56 sp99_56 78000.000000
Rwpos99_57 in99_57 sp99_57 202000.000000
Rwpos99_58 in99_58 sp99_58 78000.000000
Rwpos99_59 in99_59 sp99_59 202000.000000
Rwpos99_60 in99_60 sp99_60 78000.000000
Rwpos99_61 in99_61 sp99_61 78000.000000
Rwpos99_62 in99_62 sp99_62 78000.000000
Rwpos99_63 in99_63 sp99_63 202000.000000
Rwpos99_64 in99_64 sp99_64 202000.000000
Rwpos99_65 in99_65 sp99_65 202000.000000
Rwpos99_66 in99_66 sp99_66 202000.000000
Rwpos99_67 in99_67 sp99_67 78000.000000
Rwpos99_68 in99_68 sp99_68 78000.000000
Rwpos99_69 in99_69 sp99_69 78000.000000
Rwpos99_70 in99_70 sp99_70 202000.000000
Rwpos99_71 in99_71 sp99_71 78000.000000
Rwpos99_72 in99_72 sp99_72 202000.000000
Rwpos99_73 in99_73 sp99_73 78000.000000
Rwpos99_74 in99_74 sp99_74 78000.000000
Rwpos99_75 in99_75 sp99_75 202000.000000
Rwpos99_76 in99_76 sp99_76 202000.000000
Rwpos99_77 in99_77 sp99_77 78000.000000
Rwpos99_78 in99_78 sp99_78 78000.000000
Rwpos99_79 in99_79 sp99_79 78000.000000
Rwpos99_80 in99_80 sp99_80 78000.000000
Rwpos99_81 in99_81 sp99_81 78000.000000
Rwpos99_82 in99_82 sp99_82 78000.000000
Rwpos99_83 in99_83 sp99_83 78000.000000
Rwpos99_84 in99_84 sp99_84 202000.000000
Rwpos100_1 in100_1 sp100_1 78000.000000
Rwpos100_2 in100_2 sp100_2 78000.000000
Rwpos100_3 in100_3 sp100_3 202000.000000
Rwpos100_4 in100_4 sp100_4 202000.000000
Rwpos100_5 in100_5 sp100_5 202000.000000
Rwpos100_6 in100_6 sp100_6 78000.000000
Rwpos100_7 in100_7 sp100_7 202000.000000
Rwpos100_8 in100_8 sp100_8 202000.000000
Rwpos100_9 in100_9 sp100_9 202000.000000
Rwpos100_10 in100_10 sp100_10 202000.000000
Rwpos100_11 in100_11 sp100_11 78000.000000
Rwpos100_12 in100_12 sp100_12 78000.000000
Rwpos100_13 in100_13 sp100_13 202000.000000
Rwpos100_14 in100_14 sp100_14 202000.000000
Rwpos100_15 in100_15 sp100_15 78000.000000
Rwpos100_16 in100_16 sp100_16 78000.000000
Rwpos100_17 in100_17 sp100_17 78000.000000
Rwpos100_18 in100_18 sp100_18 78000.000000
Rwpos100_19 in100_19 sp100_19 78000.000000
Rwpos100_20 in100_20 sp100_20 78000.000000
Rwpos100_21 in100_21 sp100_21 78000.000000
Rwpos100_22 in100_22 sp100_22 202000.000000
Rwpos100_23 in100_23 sp100_23 78000.000000
Rwpos100_24 in100_24 sp100_24 202000.000000
Rwpos100_25 in100_25 sp100_25 202000.000000
Rwpos100_26 in100_26 sp100_26 202000.000000
Rwpos100_27 in100_27 sp100_27 202000.000000
Rwpos100_28 in100_28 sp100_28 78000.000000
Rwpos100_29 in100_29 sp100_29 202000.000000
Rwpos100_30 in100_30 sp100_30 78000.000000
Rwpos100_31 in100_31 sp100_31 202000.000000
Rwpos100_32 in100_32 sp100_32 78000.000000
Rwpos100_33 in100_33 sp100_33 78000.000000
Rwpos100_34 in100_34 sp100_34 202000.000000
Rwpos100_35 in100_35 sp100_35 202000.000000
Rwpos100_36 in100_36 sp100_36 202000.000000
Rwpos100_37 in100_37 sp100_37 78000.000000
Rwpos100_38 in100_38 sp100_38 78000.000000
Rwpos100_39 in100_39 sp100_39 202000.000000
Rwpos100_40 in100_40 sp100_40 78000.000000
Rwpos100_41 in100_41 sp100_41 202000.000000
Rwpos100_42 in100_42 sp100_42 78000.000000
Rwpos100_43 in100_43 sp100_43 78000.000000
Rwpos100_44 in100_44 sp100_44 202000.000000
Rwpos100_45 in100_45 sp100_45 78000.000000
Rwpos100_46 in100_46 sp100_46 78000.000000
Rwpos100_47 in100_47 sp100_47 202000.000000
Rwpos100_48 in100_48 sp100_48 202000.000000
Rwpos100_49 in100_49 sp100_49 78000.000000
Rwpos100_50 in100_50 sp100_50 202000.000000
Rwpos100_51 in100_51 sp100_51 202000.000000
Rwpos100_52 in100_52 sp100_52 78000.000000
Rwpos100_53 in100_53 sp100_53 78000.000000
Rwpos100_54 in100_54 sp100_54 78000.000000
Rwpos100_55 in100_55 sp100_55 78000.000000
Rwpos100_56 in100_56 sp100_56 78000.000000
Rwpos100_57 in100_57 sp100_57 202000.000000
Rwpos100_58 in100_58 sp100_58 78000.000000
Rwpos100_59 in100_59 sp100_59 78000.000000
Rwpos100_60 in100_60 sp100_60 202000.000000
Rwpos100_61 in100_61 sp100_61 78000.000000
Rwpos100_62 in100_62 sp100_62 202000.000000
Rwpos100_63 in100_63 sp100_63 78000.000000
Rwpos100_64 in100_64 sp100_64 78000.000000
Rwpos100_65 in100_65 sp100_65 202000.000000
Rwpos100_66 in100_66 sp100_66 202000.000000
Rwpos100_67 in100_67 sp100_67 202000.000000
Rwpos100_68 in100_68 sp100_68 78000.000000
Rwpos100_69 in100_69 sp100_69 78000.000000
Rwpos100_70 in100_70 sp100_70 202000.000000
Rwpos100_71 in100_71 sp100_71 78000.000000
Rwpos100_72 in100_72 sp100_72 202000.000000
Rwpos100_73 in100_73 sp100_73 78000.000000
Rwpos100_74 in100_74 sp100_74 202000.000000
Rwpos100_75 in100_75 sp100_75 202000.000000
Rwpos100_76 in100_76 sp100_76 202000.000000
Rwpos100_77 in100_77 sp100_77 78000.000000
Rwpos100_78 in100_78 sp100_78 202000.000000
Rwpos100_79 in100_79 sp100_79 78000.000000
Rwpos100_80 in100_80 sp100_80 78000.000000
Rwpos100_81 in100_81 sp100_81 78000.000000
Rwpos100_82 in100_82 sp100_82 202000.000000
Rwpos100_83 in100_83 sp100_83 78000.000000
Rwpos100_84 in100_84 sp100_84 78000.000000
Rwpos101_1 in101_1 sp101_1 78000.000000
Rwpos101_2 in101_2 sp101_2 78000.000000
Rwpos101_3 in101_3 sp101_3 202000.000000
Rwpos101_4 in101_4 sp101_4 202000.000000
Rwpos101_5 in101_5 sp101_5 202000.000000
Rwpos101_6 in101_6 sp101_6 78000.000000
Rwpos101_7 in101_7 sp101_7 78000.000000
Rwpos101_8 in101_8 sp101_8 78000.000000
Rwpos101_9 in101_9 sp101_9 202000.000000
Rwpos101_10 in101_10 sp101_10 78000.000000
Rwpos101_11 in101_11 sp101_11 78000.000000
Rwpos101_12 in101_12 sp101_12 202000.000000
Rwpos101_13 in101_13 sp101_13 78000.000000
Rwpos101_14 in101_14 sp101_14 78000.000000
Rwpos101_15 in101_15 sp101_15 78000.000000
Rwpos101_16 in101_16 sp101_16 202000.000000
Rwpos101_17 in101_17 sp101_17 202000.000000
Rwpos101_18 in101_18 sp101_18 202000.000000
Rwpos101_19 in101_19 sp101_19 78000.000000
Rwpos101_20 in101_20 sp101_20 78000.000000
Rwpos101_21 in101_21 sp101_21 78000.000000
Rwpos101_22 in101_22 sp101_22 202000.000000
Rwpos101_23 in101_23 sp101_23 78000.000000
Rwpos101_24 in101_24 sp101_24 78000.000000
Rwpos101_25 in101_25 sp101_25 78000.000000
Rwpos101_26 in101_26 sp101_26 202000.000000
Rwpos101_27 in101_27 sp101_27 202000.000000
Rwpos101_28 in101_28 sp101_28 78000.000000
Rwpos101_29 in101_29 sp101_29 202000.000000
Rwpos101_30 in101_30 sp101_30 78000.000000
Rwpos101_31 in101_31 sp101_31 202000.000000
Rwpos101_32 in101_32 sp101_32 202000.000000
Rwpos101_33 in101_33 sp101_33 202000.000000
Rwpos101_34 in101_34 sp101_34 78000.000000
Rwpos101_35 in101_35 sp101_35 202000.000000
Rwpos101_36 in101_36 sp101_36 78000.000000
Rwpos101_37 in101_37 sp101_37 78000.000000
Rwpos101_38 in101_38 sp101_38 78000.000000
Rwpos101_39 in101_39 sp101_39 78000.000000
Rwpos101_40 in101_40 sp101_40 202000.000000
Rwpos101_41 in101_41 sp101_41 202000.000000
Rwpos101_42 in101_42 sp101_42 78000.000000
Rwpos101_43 in101_43 sp101_43 202000.000000
Rwpos101_44 in101_44 sp101_44 78000.000000
Rwpos101_45 in101_45 sp101_45 78000.000000
Rwpos101_46 in101_46 sp101_46 78000.000000
Rwpos101_47 in101_47 sp101_47 78000.000000
Rwpos101_48 in101_48 sp101_48 78000.000000
Rwpos101_49 in101_49 sp101_49 78000.000000
Rwpos101_50 in101_50 sp101_50 78000.000000
Rwpos101_51 in101_51 sp101_51 202000.000000
Rwpos101_52 in101_52 sp101_52 78000.000000
Rwpos101_53 in101_53 sp101_53 78000.000000
Rwpos101_54 in101_54 sp101_54 202000.000000
Rwpos101_55 in101_55 sp101_55 202000.000000
Rwpos101_56 in101_56 sp101_56 78000.000000
Rwpos101_57 in101_57 sp101_57 202000.000000
Rwpos101_58 in101_58 sp101_58 78000.000000
Rwpos101_59 in101_59 sp101_59 78000.000000
Rwpos101_60 in101_60 sp101_60 78000.000000
Rwpos101_61 in101_61 sp101_61 202000.000000
Rwpos101_62 in101_62 sp101_62 202000.000000
Rwpos101_63 in101_63 sp101_63 78000.000000
Rwpos101_64 in101_64 sp101_64 202000.000000
Rwpos101_65 in101_65 sp101_65 78000.000000
Rwpos101_66 in101_66 sp101_66 202000.000000
Rwpos101_67 in101_67 sp101_67 78000.000000
Rwpos101_68 in101_68 sp101_68 202000.000000
Rwpos101_69 in101_69 sp101_69 202000.000000
Rwpos101_70 in101_70 sp101_70 202000.000000
Rwpos101_71 in101_71 sp101_71 78000.000000
Rwpos101_72 in101_72 sp101_72 202000.000000
Rwpos101_73 in101_73 sp101_73 202000.000000
Rwpos101_74 in101_74 sp101_74 202000.000000
Rwpos101_75 in101_75 sp101_75 78000.000000
Rwpos101_76 in101_76 sp101_76 78000.000000
Rwpos101_77 in101_77 sp101_77 78000.000000
Rwpos101_78 in101_78 sp101_78 202000.000000
Rwpos101_79 in101_79 sp101_79 78000.000000
Rwpos101_80 in101_80 sp101_80 202000.000000
Rwpos101_81 in101_81 sp101_81 78000.000000
Rwpos101_82 in101_82 sp101_82 78000.000000
Rwpos101_83 in101_83 sp101_83 202000.000000
Rwpos101_84 in101_84 sp101_84 78000.000000
Rwpos102_1 in102_1 sp102_1 202000.000000
Rwpos102_2 in102_2 sp102_2 78000.000000
Rwpos102_3 in102_3 sp102_3 202000.000000
Rwpos102_4 in102_4 sp102_4 78000.000000
Rwpos102_5 in102_5 sp102_5 202000.000000
Rwpos102_6 in102_6 sp102_6 78000.000000
Rwpos102_7 in102_7 sp102_7 78000.000000
Rwpos102_8 in102_8 sp102_8 78000.000000
Rwpos102_9 in102_9 sp102_9 78000.000000
Rwpos102_10 in102_10 sp102_10 78000.000000
Rwpos102_11 in102_11 sp102_11 78000.000000
Rwpos102_12 in102_12 sp102_12 202000.000000
Rwpos102_13 in102_13 sp102_13 78000.000000
Rwpos102_14 in102_14 sp102_14 202000.000000
Rwpos102_15 in102_15 sp102_15 78000.000000
Rwpos102_16 in102_16 sp102_16 202000.000000
Rwpos102_17 in102_17 sp102_17 78000.000000
Rwpos102_18 in102_18 sp102_18 202000.000000
Rwpos102_19 in102_19 sp102_19 202000.000000
Rwpos102_20 in102_20 sp102_20 202000.000000
Rwpos102_21 in102_21 sp102_21 78000.000000
Rwpos102_22 in102_22 sp102_22 78000.000000
Rwpos102_23 in102_23 sp102_23 78000.000000
Rwpos102_24 in102_24 sp102_24 78000.000000
Rwpos102_25 in102_25 sp102_25 202000.000000
Rwpos102_26 in102_26 sp102_26 202000.000000
Rwpos102_27 in102_27 sp102_27 78000.000000
Rwpos102_28 in102_28 sp102_28 202000.000000
Rwpos102_29 in102_29 sp102_29 202000.000000
Rwpos102_30 in102_30 sp102_30 78000.000000
Rwpos102_31 in102_31 sp102_31 78000.000000
Rwpos102_32 in102_32 sp102_32 202000.000000
Rwpos102_33 in102_33 sp102_33 202000.000000
Rwpos102_34 in102_34 sp102_34 202000.000000
Rwpos102_35 in102_35 sp102_35 202000.000000
Rwpos102_36 in102_36 sp102_36 78000.000000
Rwpos102_37 in102_37 sp102_37 78000.000000
Rwpos102_38 in102_38 sp102_38 202000.000000
Rwpos102_39 in102_39 sp102_39 202000.000000
Rwpos102_40 in102_40 sp102_40 202000.000000
Rwpos102_41 in102_41 sp102_41 202000.000000
Rwpos102_42 in102_42 sp102_42 202000.000000
Rwpos102_43 in102_43 sp102_43 78000.000000
Rwpos102_44 in102_44 sp102_44 78000.000000
Rwpos102_45 in102_45 sp102_45 202000.000000
Rwpos102_46 in102_46 sp102_46 202000.000000
Rwpos102_47 in102_47 sp102_47 78000.000000
Rwpos102_48 in102_48 sp102_48 202000.000000
Rwpos102_49 in102_49 sp102_49 202000.000000
Rwpos102_50 in102_50 sp102_50 202000.000000
Rwpos102_51 in102_51 sp102_51 202000.000000
Rwpos102_52 in102_52 sp102_52 78000.000000
Rwpos102_53 in102_53 sp102_53 202000.000000
Rwpos102_54 in102_54 sp102_54 202000.000000
Rwpos102_55 in102_55 sp102_55 78000.000000
Rwpos102_56 in102_56 sp102_56 78000.000000
Rwpos102_57 in102_57 sp102_57 202000.000000
Rwpos102_58 in102_58 sp102_58 78000.000000
Rwpos102_59 in102_59 sp102_59 78000.000000
Rwpos102_60 in102_60 sp102_60 78000.000000
Rwpos102_61 in102_61 sp102_61 78000.000000
Rwpos102_62 in102_62 sp102_62 78000.000000
Rwpos102_63 in102_63 sp102_63 78000.000000
Rwpos102_64 in102_64 sp102_64 78000.000000
Rwpos102_65 in102_65 sp102_65 78000.000000
Rwpos102_66 in102_66 sp102_66 78000.000000
Rwpos102_67 in102_67 sp102_67 202000.000000
Rwpos102_68 in102_68 sp102_68 78000.000000
Rwpos102_69 in102_69 sp102_69 78000.000000
Rwpos102_70 in102_70 sp102_70 78000.000000
Rwpos102_71 in102_71 sp102_71 78000.000000
Rwpos102_72 in102_72 sp102_72 78000.000000
Rwpos102_73 in102_73 sp102_73 78000.000000
Rwpos102_74 in102_74 sp102_74 78000.000000
Rwpos102_75 in102_75 sp102_75 202000.000000
Rwpos102_76 in102_76 sp102_76 78000.000000
Rwpos102_77 in102_77 sp102_77 78000.000000
Rwpos102_78 in102_78 sp102_78 78000.000000
Rwpos102_79 in102_79 sp102_79 78000.000000
Rwpos102_80 in102_80 sp102_80 202000.000000
Rwpos102_81 in102_81 sp102_81 78000.000000
Rwpos102_82 in102_82 sp102_82 78000.000000
Rwpos102_83 in102_83 sp102_83 202000.000000
Rwpos102_84 in102_84 sp102_84 202000.000000
Rwpos103_1 in103_1 sp103_1 202000.000000
Rwpos103_2 in103_2 sp103_2 202000.000000
Rwpos103_3 in103_3 sp103_3 78000.000000
Rwpos103_4 in103_4 sp103_4 202000.000000
Rwpos103_5 in103_5 sp103_5 202000.000000
Rwpos103_6 in103_6 sp103_6 202000.000000
Rwpos103_7 in103_7 sp103_7 78000.000000
Rwpos103_8 in103_8 sp103_8 78000.000000
Rwpos103_9 in103_9 sp103_9 202000.000000
Rwpos103_10 in103_10 sp103_10 78000.000000
Rwpos103_11 in103_11 sp103_11 78000.000000
Rwpos103_12 in103_12 sp103_12 202000.000000
Rwpos103_13 in103_13 sp103_13 202000.000000
Rwpos103_14 in103_14 sp103_14 78000.000000
Rwpos103_15 in103_15 sp103_15 78000.000000
Rwpos103_16 in103_16 sp103_16 202000.000000
Rwpos103_17 in103_17 sp103_17 202000.000000
Rwpos103_18 in103_18 sp103_18 202000.000000
Rwpos103_19 in103_19 sp103_19 202000.000000
Rwpos103_20 in103_20 sp103_20 78000.000000
Rwpos103_21 in103_21 sp103_21 78000.000000
Rwpos103_22 in103_22 sp103_22 202000.000000
Rwpos103_23 in103_23 sp103_23 78000.000000
Rwpos103_24 in103_24 sp103_24 202000.000000
Rwpos103_25 in103_25 sp103_25 202000.000000
Rwpos103_26 in103_26 sp103_26 78000.000000
Rwpos103_27 in103_27 sp103_27 202000.000000
Rwpos103_28 in103_28 sp103_28 78000.000000
Rwpos103_29 in103_29 sp103_29 78000.000000
Rwpos103_30 in103_30 sp103_30 78000.000000
Rwpos103_31 in103_31 sp103_31 202000.000000
Rwpos103_32 in103_32 sp103_32 78000.000000
Rwpos103_33 in103_33 sp103_33 78000.000000
Rwpos103_34 in103_34 sp103_34 78000.000000
Rwpos103_35 in103_35 sp103_35 78000.000000
Rwpos103_36 in103_36 sp103_36 202000.000000
Rwpos103_37 in103_37 sp103_37 78000.000000
Rwpos103_38 in103_38 sp103_38 78000.000000
Rwpos103_39 in103_39 sp103_39 202000.000000
Rwpos103_40 in103_40 sp103_40 78000.000000
Rwpos103_41 in103_41 sp103_41 78000.000000
Rwpos103_42 in103_42 sp103_42 78000.000000
Rwpos103_43 in103_43 sp103_43 78000.000000
Rwpos103_44 in103_44 sp103_44 202000.000000
Rwpos103_45 in103_45 sp103_45 202000.000000
Rwpos103_46 in103_46 sp103_46 78000.000000
Rwpos103_47 in103_47 sp103_47 202000.000000
Rwpos103_48 in103_48 sp103_48 78000.000000
Rwpos103_49 in103_49 sp103_49 78000.000000
Rwpos103_50 in103_50 sp103_50 202000.000000
Rwpos103_51 in103_51 sp103_51 78000.000000
Rwpos103_52 in103_52 sp103_52 78000.000000
Rwpos103_53 in103_53 sp103_53 202000.000000
Rwpos103_54 in103_54 sp103_54 78000.000000
Rwpos103_55 in103_55 sp103_55 78000.000000
Rwpos103_56 in103_56 sp103_56 78000.000000
Rwpos103_57 in103_57 sp103_57 78000.000000
Rwpos103_58 in103_58 sp103_58 202000.000000
Rwpos103_59 in103_59 sp103_59 202000.000000
Rwpos103_60 in103_60 sp103_60 202000.000000
Rwpos103_61 in103_61 sp103_61 202000.000000
Rwpos103_62 in103_62 sp103_62 78000.000000
Rwpos103_63 in103_63 sp103_63 78000.000000
Rwpos103_64 in103_64 sp103_64 78000.000000
Rwpos103_65 in103_65 sp103_65 202000.000000
Rwpos103_66 in103_66 sp103_66 202000.000000
Rwpos103_67 in103_67 sp103_67 202000.000000
Rwpos103_68 in103_68 sp103_68 202000.000000
Rwpos103_69 in103_69 sp103_69 78000.000000
Rwpos103_70 in103_70 sp103_70 78000.000000
Rwpos103_71 in103_71 sp103_71 78000.000000
Rwpos103_72 in103_72 sp103_72 78000.000000
Rwpos103_73 in103_73 sp103_73 78000.000000
Rwpos103_74 in103_74 sp103_74 202000.000000
Rwpos103_75 in103_75 sp103_75 78000.000000
Rwpos103_76 in103_76 sp103_76 78000.000000
Rwpos103_77 in103_77 sp103_77 78000.000000
Rwpos103_78 in103_78 sp103_78 202000.000000
Rwpos103_79 in103_79 sp103_79 78000.000000
Rwpos103_80 in103_80 sp103_80 78000.000000
Rwpos103_81 in103_81 sp103_81 78000.000000
Rwpos103_82 in103_82 sp103_82 202000.000000
Rwpos103_83 in103_83 sp103_83 202000.000000
Rwpos103_84 in103_84 sp103_84 78000.000000
Rwpos104_1 in104_1 sp104_1 78000.000000
Rwpos104_2 in104_2 sp104_2 78000.000000
Rwpos104_3 in104_3 sp104_3 78000.000000
Rwpos104_4 in104_4 sp104_4 78000.000000
Rwpos104_5 in104_5 sp104_5 202000.000000
Rwpos104_6 in104_6 sp104_6 202000.000000
Rwpos104_7 in104_7 sp104_7 78000.000000
Rwpos104_8 in104_8 sp104_8 78000.000000
Rwpos104_9 in104_9 sp104_9 202000.000000
Rwpos104_10 in104_10 sp104_10 202000.000000
Rwpos104_11 in104_11 sp104_11 78000.000000
Rwpos104_12 in104_12 sp104_12 202000.000000
Rwpos104_13 in104_13 sp104_13 202000.000000
Rwpos104_14 in104_14 sp104_14 78000.000000
Rwpos104_15 in104_15 sp104_15 78000.000000
Rwpos104_16 in104_16 sp104_16 78000.000000
Rwpos104_17 in104_17 sp104_17 202000.000000
Rwpos104_18 in104_18 sp104_18 202000.000000
Rwpos104_19 in104_19 sp104_19 78000.000000
Rwpos104_20 in104_20 sp104_20 78000.000000
Rwpos104_21 in104_21 sp104_21 202000.000000
Rwpos104_22 in104_22 sp104_22 78000.000000
Rwpos104_23 in104_23 sp104_23 78000.000000
Rwpos104_24 in104_24 sp104_24 202000.000000
Rwpos104_25 in104_25 sp104_25 78000.000000
Rwpos104_26 in104_26 sp104_26 202000.000000
Rwpos104_27 in104_27 sp104_27 202000.000000
Rwpos104_28 in104_28 sp104_28 202000.000000
Rwpos104_29 in104_29 sp104_29 78000.000000
Rwpos104_30 in104_30 sp104_30 78000.000000
Rwpos104_31 in104_31 sp104_31 202000.000000
Rwpos104_32 in104_32 sp104_32 78000.000000
Rwpos104_33 in104_33 sp104_33 78000.000000
Rwpos104_34 in104_34 sp104_34 78000.000000
Rwpos104_35 in104_35 sp104_35 78000.000000
Rwpos104_36 in104_36 sp104_36 202000.000000
Rwpos104_37 in104_37 sp104_37 78000.000000
Rwpos104_38 in104_38 sp104_38 78000.000000
Rwpos104_39 in104_39 sp104_39 202000.000000
Rwpos104_40 in104_40 sp104_40 78000.000000
Rwpos104_41 in104_41 sp104_41 202000.000000
Rwpos104_42 in104_42 sp104_42 78000.000000
Rwpos104_43 in104_43 sp104_43 202000.000000
Rwpos104_44 in104_44 sp104_44 202000.000000
Rwpos104_45 in104_45 sp104_45 78000.000000
Rwpos104_46 in104_46 sp104_46 78000.000000
Rwpos104_47 in104_47 sp104_47 202000.000000
Rwpos104_48 in104_48 sp104_48 202000.000000
Rwpos104_49 in104_49 sp104_49 78000.000000
Rwpos104_50 in104_50 sp104_50 78000.000000
Rwpos104_51 in104_51 sp104_51 202000.000000
Rwpos104_52 in104_52 sp104_52 78000.000000
Rwpos104_53 in104_53 sp104_53 78000.000000
Rwpos104_54 in104_54 sp104_54 202000.000000
Rwpos104_55 in104_55 sp104_55 78000.000000
Rwpos104_56 in104_56 sp104_56 202000.000000
Rwpos104_57 in104_57 sp104_57 78000.000000
Rwpos104_58 in104_58 sp104_58 78000.000000
Rwpos104_59 in104_59 sp104_59 78000.000000
Rwpos104_60 in104_60 sp104_60 202000.000000
Rwpos104_61 in104_61 sp104_61 78000.000000
Rwpos104_62 in104_62 sp104_62 202000.000000
Rwpos104_63 in104_63 sp104_63 202000.000000
Rwpos104_64 in104_64 sp104_64 202000.000000
Rwpos104_65 in104_65 sp104_65 202000.000000
Rwpos104_66 in104_66 sp104_66 78000.000000
Rwpos104_67 in104_67 sp104_67 202000.000000
Rwpos104_68 in104_68 sp104_68 202000.000000
Rwpos104_69 in104_69 sp104_69 202000.000000
Rwpos104_70 in104_70 sp104_70 78000.000000
Rwpos104_71 in104_71 sp104_71 78000.000000
Rwpos104_72 in104_72 sp104_72 202000.000000
Rwpos104_73 in104_73 sp104_73 78000.000000
Rwpos104_74 in104_74 sp104_74 78000.000000
Rwpos104_75 in104_75 sp104_75 78000.000000
Rwpos104_76 in104_76 sp104_76 78000.000000
Rwpos104_77 in104_77 sp104_77 202000.000000
Rwpos104_78 in104_78 sp104_78 202000.000000
Rwpos104_79 in104_79 sp104_79 202000.000000
Rwpos104_80 in104_80 sp104_80 202000.000000
Rwpos104_81 in104_81 sp104_81 202000.000000
Rwpos104_82 in104_82 sp104_82 202000.000000
Rwpos104_83 in104_83 sp104_83 78000.000000
Rwpos104_84 in104_84 sp104_84 78000.000000
Rwpos105_1 in105_1 sp105_1 202000.000000
Rwpos105_2 in105_2 sp105_2 78000.000000
Rwpos105_3 in105_3 sp105_3 78000.000000
Rwpos105_4 in105_4 sp105_4 78000.000000
Rwpos105_5 in105_5 sp105_5 78000.000000
Rwpos105_6 in105_6 sp105_6 202000.000000
Rwpos105_7 in105_7 sp105_7 202000.000000
Rwpos105_8 in105_8 sp105_8 78000.000000
Rwpos105_9 in105_9 sp105_9 78000.000000
Rwpos105_10 in105_10 sp105_10 78000.000000
Rwpos105_11 in105_11 sp105_11 202000.000000
Rwpos105_12 in105_12 sp105_12 78000.000000
Rwpos105_13 in105_13 sp105_13 202000.000000
Rwpos105_14 in105_14 sp105_14 202000.000000
Rwpos105_15 in105_15 sp105_15 202000.000000
Rwpos105_16 in105_16 sp105_16 78000.000000
Rwpos105_17 in105_17 sp105_17 202000.000000
Rwpos105_18 in105_18 sp105_18 78000.000000
Rwpos105_19 in105_19 sp105_19 78000.000000
Rwpos105_20 in105_20 sp105_20 78000.000000
Rwpos105_21 in105_21 sp105_21 202000.000000
Rwpos105_22 in105_22 sp105_22 202000.000000
Rwpos105_23 in105_23 sp105_23 202000.000000
Rwpos105_24 in105_24 sp105_24 202000.000000
Rwpos105_25 in105_25 sp105_25 78000.000000
Rwpos105_26 in105_26 sp105_26 202000.000000
Rwpos105_27 in105_27 sp105_27 78000.000000
Rwpos105_28 in105_28 sp105_28 202000.000000
Rwpos105_29 in105_29 sp105_29 78000.000000
Rwpos105_30 in105_30 sp105_30 202000.000000
Rwpos105_31 in105_31 sp105_31 202000.000000
Rwpos105_32 in105_32 sp105_32 78000.000000
Rwpos105_33 in105_33 sp105_33 202000.000000
Rwpos105_34 in105_34 sp105_34 78000.000000
Rwpos105_35 in105_35 sp105_35 78000.000000
Rwpos105_36 in105_36 sp105_36 78000.000000
Rwpos105_37 in105_37 sp105_37 78000.000000
Rwpos105_38 in105_38 sp105_38 78000.000000
Rwpos105_39 in105_39 sp105_39 78000.000000
Rwpos105_40 in105_40 sp105_40 78000.000000
Rwpos105_41 in105_41 sp105_41 202000.000000
Rwpos105_42 in105_42 sp105_42 78000.000000
Rwpos105_43 in105_43 sp105_43 202000.000000
Rwpos105_44 in105_44 sp105_44 202000.000000
Rwpos105_45 in105_45 sp105_45 78000.000000
Rwpos105_46 in105_46 sp105_46 202000.000000
Rwpos105_47 in105_47 sp105_47 202000.000000
Rwpos105_48 in105_48 sp105_48 202000.000000
Rwpos105_49 in105_49 sp105_49 78000.000000
Rwpos105_50 in105_50 sp105_50 78000.000000
Rwpos105_51 in105_51 sp105_51 78000.000000
Rwpos105_52 in105_52 sp105_52 78000.000000
Rwpos105_53 in105_53 sp105_53 78000.000000
Rwpos105_54 in105_54 sp105_54 78000.000000
Rwpos105_55 in105_55 sp105_55 78000.000000
Rwpos105_56 in105_56 sp105_56 78000.000000
Rwpos105_57 in105_57 sp105_57 202000.000000
Rwpos105_58 in105_58 sp105_58 78000.000000
Rwpos105_59 in105_59 sp105_59 78000.000000
Rwpos105_60 in105_60 sp105_60 202000.000000
Rwpos105_61 in105_61 sp105_61 78000.000000
Rwpos105_62 in105_62 sp105_62 202000.000000
Rwpos105_63 in105_63 sp105_63 78000.000000
Rwpos105_64 in105_64 sp105_64 78000.000000
Rwpos105_65 in105_65 sp105_65 78000.000000
Rwpos105_66 in105_66 sp105_66 78000.000000
Rwpos105_67 in105_67 sp105_67 78000.000000
Rwpos105_68 in105_68 sp105_68 202000.000000
Rwpos105_69 in105_69 sp105_69 78000.000000
Rwpos105_70 in105_70 sp105_70 78000.000000
Rwpos105_71 in105_71 sp105_71 78000.000000
Rwpos105_72 in105_72 sp105_72 202000.000000
Rwpos105_73 in105_73 sp105_73 202000.000000
Rwpos105_74 in105_74 sp105_74 78000.000000
Rwpos105_75 in105_75 sp105_75 78000.000000
Rwpos105_76 in105_76 sp105_76 78000.000000
Rwpos105_77 in105_77 sp105_77 78000.000000
Rwpos105_78 in105_78 sp105_78 202000.000000
Rwpos105_79 in105_79 sp105_79 78000.000000
Rwpos105_80 in105_80 sp105_80 78000.000000
Rwpos105_81 in105_81 sp105_81 202000.000000
Rwpos105_82 in105_82 sp105_82 78000.000000
Rwpos105_83 in105_83 sp105_83 78000.000000
Rwpos105_84 in105_84 sp105_84 78000.000000
Rwpos106_1 in106_1 sp106_1 78000.000000
Rwpos106_2 in106_2 sp106_2 78000.000000
Rwpos106_3 in106_3 sp106_3 202000.000000
Rwpos106_4 in106_4 sp106_4 78000.000000
Rwpos106_5 in106_5 sp106_5 202000.000000
Rwpos106_6 in106_6 sp106_6 78000.000000
Rwpos106_7 in106_7 sp106_7 78000.000000
Rwpos106_8 in106_8 sp106_8 202000.000000
Rwpos106_9 in106_9 sp106_9 202000.000000
Rwpos106_10 in106_10 sp106_10 78000.000000
Rwpos106_11 in106_11 sp106_11 202000.000000
Rwpos106_12 in106_12 sp106_12 78000.000000
Rwpos106_13 in106_13 sp106_13 202000.000000
Rwpos106_14 in106_14 sp106_14 78000.000000
Rwpos106_15 in106_15 sp106_15 202000.000000
Rwpos106_16 in106_16 sp106_16 78000.000000
Rwpos106_17 in106_17 sp106_17 78000.000000
Rwpos106_18 in106_18 sp106_18 202000.000000
Rwpos106_19 in106_19 sp106_19 78000.000000
Rwpos106_20 in106_20 sp106_20 202000.000000
Rwpos106_21 in106_21 sp106_21 202000.000000
Rwpos106_22 in106_22 sp106_22 78000.000000
Rwpos106_23 in106_23 sp106_23 202000.000000
Rwpos106_24 in106_24 sp106_24 78000.000000
Rwpos106_25 in106_25 sp106_25 202000.000000
Rwpos106_26 in106_26 sp106_26 202000.000000
Rwpos106_27 in106_27 sp106_27 78000.000000
Rwpos106_28 in106_28 sp106_28 78000.000000
Rwpos106_29 in106_29 sp106_29 202000.000000
Rwpos106_30 in106_30 sp106_30 78000.000000
Rwpos106_31 in106_31 sp106_31 78000.000000
Rwpos106_32 in106_32 sp106_32 78000.000000
Rwpos106_33 in106_33 sp106_33 202000.000000
Rwpos106_34 in106_34 sp106_34 202000.000000
Rwpos106_35 in106_35 sp106_35 202000.000000
Rwpos106_36 in106_36 sp106_36 78000.000000
Rwpos106_37 in106_37 sp106_37 78000.000000
Rwpos106_38 in106_38 sp106_38 78000.000000
Rwpos106_39 in106_39 sp106_39 202000.000000
Rwpos106_40 in106_40 sp106_40 78000.000000
Rwpos106_41 in106_41 sp106_41 202000.000000
Rwpos106_42 in106_42 sp106_42 78000.000000
Rwpos106_43 in106_43 sp106_43 202000.000000
Rwpos106_44 in106_44 sp106_44 78000.000000
Rwpos106_45 in106_45 sp106_45 78000.000000
Rwpos106_46 in106_46 sp106_46 78000.000000
Rwpos106_47 in106_47 sp106_47 78000.000000
Rwpos106_48 in106_48 sp106_48 202000.000000
Rwpos106_49 in106_49 sp106_49 78000.000000
Rwpos106_50 in106_50 sp106_50 78000.000000
Rwpos106_51 in106_51 sp106_51 78000.000000
Rwpos106_52 in106_52 sp106_52 78000.000000
Rwpos106_53 in106_53 sp106_53 202000.000000
Rwpos106_54 in106_54 sp106_54 78000.000000
Rwpos106_55 in106_55 sp106_55 202000.000000
Rwpos106_56 in106_56 sp106_56 202000.000000
Rwpos106_57 in106_57 sp106_57 78000.000000
Rwpos106_58 in106_58 sp106_58 78000.000000
Rwpos106_59 in106_59 sp106_59 202000.000000
Rwpos106_60 in106_60 sp106_60 78000.000000
Rwpos106_61 in106_61 sp106_61 202000.000000
Rwpos106_62 in106_62 sp106_62 78000.000000
Rwpos106_63 in106_63 sp106_63 202000.000000
Rwpos106_64 in106_64 sp106_64 202000.000000
Rwpos106_65 in106_65 sp106_65 202000.000000
Rwpos106_66 in106_66 sp106_66 78000.000000
Rwpos106_67 in106_67 sp106_67 78000.000000
Rwpos106_68 in106_68 sp106_68 78000.000000
Rwpos106_69 in106_69 sp106_69 202000.000000
Rwpos106_70 in106_70 sp106_70 78000.000000
Rwpos106_71 in106_71 sp106_71 202000.000000
Rwpos106_72 in106_72 sp106_72 78000.000000
Rwpos106_73 in106_73 sp106_73 202000.000000
Rwpos106_74 in106_74 sp106_74 202000.000000
Rwpos106_75 in106_75 sp106_75 202000.000000
Rwpos106_76 in106_76 sp106_76 78000.000000
Rwpos106_77 in106_77 sp106_77 202000.000000
Rwpos106_78 in106_78 sp106_78 78000.000000
Rwpos106_79 in106_79 sp106_79 202000.000000
Rwpos106_80 in106_80 sp106_80 202000.000000
Rwpos106_81 in106_81 sp106_81 202000.000000
Rwpos106_82 in106_82 sp106_82 202000.000000
Rwpos106_83 in106_83 sp106_83 202000.000000
Rwpos106_84 in106_84 sp106_84 202000.000000
Rwpos107_1 in107_1 sp107_1 78000.000000
Rwpos107_2 in107_2 sp107_2 78000.000000
Rwpos107_3 in107_3 sp107_3 78000.000000
Rwpos107_4 in107_4 sp107_4 78000.000000
Rwpos107_5 in107_5 sp107_5 78000.000000
Rwpos107_6 in107_6 sp107_6 78000.000000
Rwpos107_7 in107_7 sp107_7 202000.000000
Rwpos107_8 in107_8 sp107_8 202000.000000
Rwpos107_9 in107_9 sp107_9 78000.000000
Rwpos107_10 in107_10 sp107_10 202000.000000
Rwpos107_11 in107_11 sp107_11 202000.000000
Rwpos107_12 in107_12 sp107_12 202000.000000
Rwpos107_13 in107_13 sp107_13 78000.000000
Rwpos107_14 in107_14 sp107_14 78000.000000
Rwpos107_15 in107_15 sp107_15 78000.000000
Rwpos107_16 in107_16 sp107_16 78000.000000
Rwpos107_17 in107_17 sp107_17 78000.000000
Rwpos107_18 in107_18 sp107_18 202000.000000
Rwpos107_19 in107_19 sp107_19 78000.000000
Rwpos107_20 in107_20 sp107_20 202000.000000
Rwpos107_21 in107_21 sp107_21 78000.000000
Rwpos107_22 in107_22 sp107_22 78000.000000
Rwpos107_23 in107_23 sp107_23 202000.000000
Rwpos107_24 in107_24 sp107_24 78000.000000
Rwpos107_25 in107_25 sp107_25 78000.000000
Rwpos107_26 in107_26 sp107_26 78000.000000
Rwpos107_27 in107_27 sp107_27 78000.000000
Rwpos107_28 in107_28 sp107_28 78000.000000
Rwpos107_29 in107_29 sp107_29 202000.000000
Rwpos107_30 in107_30 sp107_30 78000.000000
Rwpos107_31 in107_31 sp107_31 78000.000000
Rwpos107_32 in107_32 sp107_32 202000.000000
Rwpos107_33 in107_33 sp107_33 78000.000000
Rwpos107_34 in107_34 sp107_34 202000.000000
Rwpos107_35 in107_35 sp107_35 78000.000000
Rwpos107_36 in107_36 sp107_36 202000.000000
Rwpos107_37 in107_37 sp107_37 202000.000000
Rwpos107_38 in107_38 sp107_38 78000.000000
Rwpos107_39 in107_39 sp107_39 202000.000000
Rwpos107_40 in107_40 sp107_40 202000.000000
Rwpos107_41 in107_41 sp107_41 78000.000000
Rwpos107_42 in107_42 sp107_42 78000.000000
Rwpos107_43 in107_43 sp107_43 78000.000000
Rwpos107_44 in107_44 sp107_44 78000.000000
Rwpos107_45 in107_45 sp107_45 78000.000000
Rwpos107_46 in107_46 sp107_46 202000.000000
Rwpos107_47 in107_47 sp107_47 78000.000000
Rwpos107_48 in107_48 sp107_48 202000.000000
Rwpos107_49 in107_49 sp107_49 202000.000000
Rwpos107_50 in107_50 sp107_50 78000.000000
Rwpos107_51 in107_51 sp107_51 78000.000000
Rwpos107_52 in107_52 sp107_52 202000.000000
Rwpos107_53 in107_53 sp107_53 202000.000000
Rwpos107_54 in107_54 sp107_54 78000.000000
Rwpos107_55 in107_55 sp107_55 202000.000000
Rwpos107_56 in107_56 sp107_56 202000.000000
Rwpos107_57 in107_57 sp107_57 202000.000000
Rwpos107_58 in107_58 sp107_58 202000.000000
Rwpos107_59 in107_59 sp107_59 78000.000000
Rwpos107_60 in107_60 sp107_60 78000.000000
Rwpos107_61 in107_61 sp107_61 202000.000000
Rwpos107_62 in107_62 sp107_62 78000.000000
Rwpos107_63 in107_63 sp107_63 202000.000000
Rwpos107_64 in107_64 sp107_64 202000.000000
Rwpos107_65 in107_65 sp107_65 202000.000000
Rwpos107_66 in107_66 sp107_66 202000.000000
Rwpos107_67 in107_67 sp107_67 78000.000000
Rwpos107_68 in107_68 sp107_68 202000.000000
Rwpos107_69 in107_69 sp107_69 202000.000000
Rwpos107_70 in107_70 sp107_70 78000.000000
Rwpos107_71 in107_71 sp107_71 202000.000000
Rwpos107_72 in107_72 sp107_72 78000.000000
Rwpos107_73 in107_73 sp107_73 202000.000000
Rwpos107_74 in107_74 sp107_74 78000.000000
Rwpos107_75 in107_75 sp107_75 202000.000000
Rwpos107_76 in107_76 sp107_76 202000.000000
Rwpos107_77 in107_77 sp107_77 202000.000000
Rwpos107_78 in107_78 sp107_78 78000.000000
Rwpos107_79 in107_79 sp107_79 202000.000000
Rwpos107_80 in107_80 sp107_80 202000.000000
Rwpos107_81 in107_81 sp107_81 78000.000000
Rwpos107_82 in107_82 sp107_82 202000.000000
Rwpos107_83 in107_83 sp107_83 202000.000000
Rwpos107_84 in107_84 sp107_84 78000.000000
Rwpos108_1 in108_1 sp108_1 78000.000000
Rwpos108_2 in108_2 sp108_2 78000.000000
Rwpos108_3 in108_3 sp108_3 78000.000000
Rwpos108_4 in108_4 sp108_4 78000.000000
Rwpos108_5 in108_5 sp108_5 78000.000000
Rwpos108_6 in108_6 sp108_6 78000.000000
Rwpos108_7 in108_7 sp108_7 78000.000000
Rwpos108_8 in108_8 sp108_8 78000.000000
Rwpos108_9 in108_9 sp108_9 78000.000000
Rwpos108_10 in108_10 sp108_10 202000.000000
Rwpos108_11 in108_11 sp108_11 78000.000000
Rwpos108_12 in108_12 sp108_12 78000.000000
Rwpos108_13 in108_13 sp108_13 78000.000000
Rwpos108_14 in108_14 sp108_14 78000.000000
Rwpos108_15 in108_15 sp108_15 202000.000000
Rwpos108_16 in108_16 sp108_16 202000.000000
Rwpos108_17 in108_17 sp108_17 78000.000000
Rwpos108_18 in108_18 sp108_18 202000.000000
Rwpos108_19 in108_19 sp108_19 202000.000000
Rwpos108_20 in108_20 sp108_20 202000.000000
Rwpos108_21 in108_21 sp108_21 78000.000000
Rwpos108_22 in108_22 sp108_22 78000.000000
Rwpos108_23 in108_23 sp108_23 202000.000000
Rwpos108_24 in108_24 sp108_24 78000.000000
Rwpos108_25 in108_25 sp108_25 202000.000000
Rwpos108_26 in108_26 sp108_26 202000.000000
Rwpos108_27 in108_27 sp108_27 78000.000000
Rwpos108_28 in108_28 sp108_28 202000.000000
Rwpos108_29 in108_29 sp108_29 78000.000000
Rwpos108_30 in108_30 sp108_30 78000.000000
Rwpos108_31 in108_31 sp108_31 78000.000000
Rwpos108_32 in108_32 sp108_32 78000.000000
Rwpos108_33 in108_33 sp108_33 202000.000000
Rwpos108_34 in108_34 sp108_34 78000.000000
Rwpos108_35 in108_35 sp108_35 78000.000000
Rwpos108_36 in108_36 sp108_36 78000.000000
Rwpos108_37 in108_37 sp108_37 202000.000000
Rwpos108_38 in108_38 sp108_38 202000.000000
Rwpos108_39 in108_39 sp108_39 202000.000000
Rwpos108_40 in108_40 sp108_40 202000.000000
Rwpos108_41 in108_41 sp108_41 202000.000000
Rwpos108_42 in108_42 sp108_42 78000.000000
Rwpos108_43 in108_43 sp108_43 202000.000000
Rwpos108_44 in108_44 sp108_44 78000.000000
Rwpos108_45 in108_45 sp108_45 202000.000000
Rwpos108_46 in108_46 sp108_46 78000.000000
Rwpos108_47 in108_47 sp108_47 78000.000000
Rwpos108_48 in108_48 sp108_48 78000.000000
Rwpos108_49 in108_49 sp108_49 202000.000000
Rwpos108_50 in108_50 sp108_50 78000.000000
Rwpos108_51 in108_51 sp108_51 202000.000000
Rwpos108_52 in108_52 sp108_52 78000.000000
Rwpos108_53 in108_53 sp108_53 202000.000000
Rwpos108_54 in108_54 sp108_54 78000.000000
Rwpos108_55 in108_55 sp108_55 202000.000000
Rwpos108_56 in108_56 sp108_56 202000.000000
Rwpos108_57 in108_57 sp108_57 78000.000000
Rwpos108_58 in108_58 sp108_58 78000.000000
Rwpos108_59 in108_59 sp108_59 78000.000000
Rwpos108_60 in108_60 sp108_60 78000.000000
Rwpos108_61 in108_61 sp108_61 78000.000000
Rwpos108_62 in108_62 sp108_62 78000.000000
Rwpos108_63 in108_63 sp108_63 202000.000000
Rwpos108_64 in108_64 sp108_64 202000.000000
Rwpos108_65 in108_65 sp108_65 202000.000000
Rwpos108_66 in108_66 sp108_66 78000.000000
Rwpos108_67 in108_67 sp108_67 78000.000000
Rwpos108_68 in108_68 sp108_68 78000.000000
Rwpos108_69 in108_69 sp108_69 78000.000000
Rwpos108_70 in108_70 sp108_70 202000.000000
Rwpos108_71 in108_71 sp108_71 202000.000000
Rwpos108_72 in108_72 sp108_72 78000.000000
Rwpos108_73 in108_73 sp108_73 78000.000000
Rwpos108_74 in108_74 sp108_74 78000.000000
Rwpos108_75 in108_75 sp108_75 202000.000000
Rwpos108_76 in108_76 sp108_76 78000.000000
Rwpos108_77 in108_77 sp108_77 202000.000000
Rwpos108_78 in108_78 sp108_78 78000.000000
Rwpos108_79 in108_79 sp108_79 78000.000000
Rwpos108_80 in108_80 sp108_80 202000.000000
Rwpos108_81 in108_81 sp108_81 78000.000000
Rwpos108_82 in108_82 sp108_82 78000.000000
Rwpos108_83 in108_83 sp108_83 78000.000000
Rwpos108_84 in108_84 sp108_84 202000.000000
Rwpos109_1 in109_1 sp109_1 202000.000000
Rwpos109_2 in109_2 sp109_2 202000.000000
Rwpos109_3 in109_3 sp109_3 202000.000000
Rwpos109_4 in109_4 sp109_4 202000.000000
Rwpos109_5 in109_5 sp109_5 202000.000000
Rwpos109_6 in109_6 sp109_6 202000.000000
Rwpos109_7 in109_7 sp109_7 78000.000000
Rwpos109_8 in109_8 sp109_8 202000.000000
Rwpos109_9 in109_9 sp109_9 78000.000000
Rwpos109_10 in109_10 sp109_10 78000.000000
Rwpos109_11 in109_11 sp109_11 78000.000000
Rwpos109_12 in109_12 sp109_12 202000.000000
Rwpos109_13 in109_13 sp109_13 202000.000000
Rwpos109_14 in109_14 sp109_14 202000.000000
Rwpos109_15 in109_15 sp109_15 78000.000000
Rwpos109_16 in109_16 sp109_16 202000.000000
Rwpos109_17 in109_17 sp109_17 78000.000000
Rwpos109_18 in109_18 sp109_18 202000.000000
Rwpos109_19 in109_19 sp109_19 202000.000000
Rwpos109_20 in109_20 sp109_20 78000.000000
Rwpos109_21 in109_21 sp109_21 202000.000000
Rwpos109_22 in109_22 sp109_22 202000.000000
Rwpos109_23 in109_23 sp109_23 78000.000000
Rwpos109_24 in109_24 sp109_24 78000.000000
Rwpos109_25 in109_25 sp109_25 202000.000000
Rwpos109_26 in109_26 sp109_26 78000.000000
Rwpos109_27 in109_27 sp109_27 202000.000000
Rwpos109_28 in109_28 sp109_28 78000.000000
Rwpos109_29 in109_29 sp109_29 78000.000000
Rwpos109_30 in109_30 sp109_30 202000.000000
Rwpos109_31 in109_31 sp109_31 202000.000000
Rwpos109_32 in109_32 sp109_32 78000.000000
Rwpos109_33 in109_33 sp109_33 78000.000000
Rwpos109_34 in109_34 sp109_34 78000.000000
Rwpos109_35 in109_35 sp109_35 202000.000000
Rwpos109_36 in109_36 sp109_36 78000.000000
Rwpos109_37 in109_37 sp109_37 78000.000000
Rwpos109_38 in109_38 sp109_38 202000.000000
Rwpos109_39 in109_39 sp109_39 202000.000000
Rwpos109_40 in109_40 sp109_40 78000.000000
Rwpos109_41 in109_41 sp109_41 202000.000000
Rwpos109_42 in109_42 sp109_42 202000.000000
Rwpos109_43 in109_43 sp109_43 202000.000000
Rwpos109_44 in109_44 sp109_44 202000.000000
Rwpos109_45 in109_45 sp109_45 202000.000000
Rwpos109_46 in109_46 sp109_46 78000.000000
Rwpos109_47 in109_47 sp109_47 202000.000000
Rwpos109_48 in109_48 sp109_48 202000.000000
Rwpos109_49 in109_49 sp109_49 202000.000000
Rwpos109_50 in109_50 sp109_50 78000.000000
Rwpos109_51 in109_51 sp109_51 78000.000000
Rwpos109_52 in109_52 sp109_52 78000.000000
Rwpos109_53 in109_53 sp109_53 78000.000000
Rwpos109_54 in109_54 sp109_54 78000.000000
Rwpos109_55 in109_55 sp109_55 202000.000000
Rwpos109_56 in109_56 sp109_56 78000.000000
Rwpos109_57 in109_57 sp109_57 78000.000000
Rwpos109_58 in109_58 sp109_58 78000.000000
Rwpos109_59 in109_59 sp109_59 202000.000000
Rwpos109_60 in109_60 sp109_60 78000.000000
Rwpos109_61 in109_61 sp109_61 202000.000000
Rwpos109_62 in109_62 sp109_62 78000.000000
Rwpos109_63 in109_63 sp109_63 78000.000000
Rwpos109_64 in109_64 sp109_64 202000.000000
Rwpos109_65 in109_65 sp109_65 78000.000000
Rwpos109_66 in109_66 sp109_66 78000.000000
Rwpos109_67 in109_67 sp109_67 202000.000000
Rwpos109_68 in109_68 sp109_68 78000.000000
Rwpos109_69 in109_69 sp109_69 78000.000000
Rwpos109_70 in109_70 sp109_70 202000.000000
Rwpos109_71 in109_71 sp109_71 78000.000000
Rwpos109_72 in109_72 sp109_72 202000.000000
Rwpos109_73 in109_73 sp109_73 78000.000000
Rwpos109_74 in109_74 sp109_74 202000.000000
Rwpos109_75 in109_75 sp109_75 202000.000000
Rwpos109_76 in109_76 sp109_76 202000.000000
Rwpos109_77 in109_77 sp109_77 78000.000000
Rwpos109_78 in109_78 sp109_78 78000.000000
Rwpos109_79 in109_79 sp109_79 78000.000000
Rwpos109_80 in109_80 sp109_80 78000.000000
Rwpos109_81 in109_81 sp109_81 78000.000000
Rwpos109_82 in109_82 sp109_82 78000.000000
Rwpos109_83 in109_83 sp109_83 202000.000000
Rwpos109_84 in109_84 sp109_84 78000.000000
Rwpos110_1 in110_1 sp110_1 78000.000000
Rwpos110_2 in110_2 sp110_2 202000.000000
Rwpos110_3 in110_3 sp110_3 78000.000000
Rwpos110_4 in110_4 sp110_4 78000.000000
Rwpos110_5 in110_5 sp110_5 78000.000000
Rwpos110_6 in110_6 sp110_6 202000.000000
Rwpos110_7 in110_7 sp110_7 202000.000000
Rwpos110_8 in110_8 sp110_8 202000.000000
Rwpos110_9 in110_9 sp110_9 78000.000000
Rwpos110_10 in110_10 sp110_10 78000.000000
Rwpos110_11 in110_11 sp110_11 78000.000000
Rwpos110_12 in110_12 sp110_12 202000.000000
Rwpos110_13 in110_13 sp110_13 78000.000000
Rwpos110_14 in110_14 sp110_14 202000.000000
Rwpos110_15 in110_15 sp110_15 202000.000000
Rwpos110_16 in110_16 sp110_16 202000.000000
Rwpos110_17 in110_17 sp110_17 78000.000000
Rwpos110_18 in110_18 sp110_18 78000.000000
Rwpos110_19 in110_19 sp110_19 202000.000000
Rwpos110_20 in110_20 sp110_20 202000.000000
Rwpos110_21 in110_21 sp110_21 78000.000000
Rwpos110_22 in110_22 sp110_22 78000.000000
Rwpos110_23 in110_23 sp110_23 78000.000000
Rwpos110_24 in110_24 sp110_24 78000.000000
Rwpos110_25 in110_25 sp110_25 202000.000000
Rwpos110_26 in110_26 sp110_26 78000.000000
Rwpos110_27 in110_27 sp110_27 202000.000000
Rwpos110_28 in110_28 sp110_28 202000.000000
Rwpos110_29 in110_29 sp110_29 202000.000000
Rwpos110_30 in110_30 sp110_30 78000.000000
Rwpos110_31 in110_31 sp110_31 78000.000000
Rwpos110_32 in110_32 sp110_32 202000.000000
Rwpos110_33 in110_33 sp110_33 78000.000000
Rwpos110_34 in110_34 sp110_34 202000.000000
Rwpos110_35 in110_35 sp110_35 78000.000000
Rwpos110_36 in110_36 sp110_36 202000.000000
Rwpos110_37 in110_37 sp110_37 202000.000000
Rwpos110_38 in110_38 sp110_38 202000.000000
Rwpos110_39 in110_39 sp110_39 202000.000000
Rwpos110_40 in110_40 sp110_40 202000.000000
Rwpos110_41 in110_41 sp110_41 202000.000000
Rwpos110_42 in110_42 sp110_42 202000.000000
Rwpos110_43 in110_43 sp110_43 78000.000000
Rwpos110_44 in110_44 sp110_44 78000.000000
Rwpos110_45 in110_45 sp110_45 202000.000000
Rwpos110_46 in110_46 sp110_46 202000.000000
Rwpos110_47 in110_47 sp110_47 78000.000000
Rwpos110_48 in110_48 sp110_48 78000.000000
Rwpos110_49 in110_49 sp110_49 202000.000000
Rwpos110_50 in110_50 sp110_50 202000.000000
Rwpos110_51 in110_51 sp110_51 202000.000000
Rwpos110_52 in110_52 sp110_52 202000.000000
Rwpos110_53 in110_53 sp110_53 78000.000000
Rwpos110_54 in110_54 sp110_54 78000.000000
Rwpos110_55 in110_55 sp110_55 78000.000000
Rwpos110_56 in110_56 sp110_56 78000.000000
Rwpos110_57 in110_57 sp110_57 78000.000000
Rwpos110_58 in110_58 sp110_58 78000.000000
Rwpos110_59 in110_59 sp110_59 78000.000000
Rwpos110_60 in110_60 sp110_60 78000.000000
Rwpos110_61 in110_61 sp110_61 78000.000000
Rwpos110_62 in110_62 sp110_62 78000.000000
Rwpos110_63 in110_63 sp110_63 202000.000000
Rwpos110_64 in110_64 sp110_64 202000.000000
Rwpos110_65 in110_65 sp110_65 78000.000000
Rwpos110_66 in110_66 sp110_66 78000.000000
Rwpos110_67 in110_67 sp110_67 202000.000000
Rwpos110_68 in110_68 sp110_68 202000.000000
Rwpos110_69 in110_69 sp110_69 202000.000000
Rwpos110_70 in110_70 sp110_70 78000.000000
Rwpos110_71 in110_71 sp110_71 78000.000000
Rwpos110_72 in110_72 sp110_72 78000.000000
Rwpos110_73 in110_73 sp110_73 78000.000000
Rwpos110_74 in110_74 sp110_74 202000.000000
Rwpos110_75 in110_75 sp110_75 78000.000000
Rwpos110_76 in110_76 sp110_76 202000.000000
Rwpos110_77 in110_77 sp110_77 78000.000000
Rwpos110_78 in110_78 sp110_78 78000.000000
Rwpos110_79 in110_79 sp110_79 202000.000000
Rwpos110_80 in110_80 sp110_80 78000.000000
Rwpos110_81 in110_81 sp110_81 78000.000000
Rwpos110_82 in110_82 sp110_82 78000.000000
Rwpos110_83 in110_83 sp110_83 78000.000000
Rwpos110_84 in110_84 sp110_84 78000.000000
Rwpos111_1 in111_1 sp111_1 78000.000000
Rwpos111_2 in111_2 sp111_2 78000.000000
Rwpos111_3 in111_3 sp111_3 78000.000000
Rwpos111_4 in111_4 sp111_4 202000.000000
Rwpos111_5 in111_5 sp111_5 202000.000000
Rwpos111_6 in111_6 sp111_6 202000.000000
Rwpos111_7 in111_7 sp111_7 78000.000000
Rwpos111_8 in111_8 sp111_8 78000.000000
Rwpos111_9 in111_9 sp111_9 202000.000000
Rwpos111_10 in111_10 sp111_10 202000.000000
Rwpos111_11 in111_11 sp111_11 78000.000000
Rwpos111_12 in111_12 sp111_12 202000.000000
Rwpos111_13 in111_13 sp111_13 202000.000000
Rwpos111_14 in111_14 sp111_14 78000.000000
Rwpos111_15 in111_15 sp111_15 202000.000000
Rwpos111_16 in111_16 sp111_16 202000.000000
Rwpos111_17 in111_17 sp111_17 78000.000000
Rwpos111_18 in111_18 sp111_18 202000.000000
Rwpos111_19 in111_19 sp111_19 202000.000000
Rwpos111_20 in111_20 sp111_20 202000.000000
Rwpos111_21 in111_21 sp111_21 202000.000000
Rwpos111_22 in111_22 sp111_22 202000.000000
Rwpos111_23 in111_23 sp111_23 78000.000000
Rwpos111_24 in111_24 sp111_24 202000.000000
Rwpos111_25 in111_25 sp111_25 78000.000000
Rwpos111_26 in111_26 sp111_26 202000.000000
Rwpos111_27 in111_27 sp111_27 202000.000000
Rwpos111_28 in111_28 sp111_28 202000.000000
Rwpos111_29 in111_29 sp111_29 202000.000000
Rwpos111_30 in111_30 sp111_30 78000.000000
Rwpos111_31 in111_31 sp111_31 78000.000000
Rwpos111_32 in111_32 sp111_32 78000.000000
Rwpos111_33 in111_33 sp111_33 202000.000000
Rwpos111_34 in111_34 sp111_34 78000.000000
Rwpos111_35 in111_35 sp111_35 202000.000000
Rwpos111_36 in111_36 sp111_36 202000.000000
Rwpos111_37 in111_37 sp111_37 78000.000000
Rwpos111_38 in111_38 sp111_38 202000.000000
Rwpos111_39 in111_39 sp111_39 202000.000000
Rwpos111_40 in111_40 sp111_40 202000.000000
Rwpos111_41 in111_41 sp111_41 202000.000000
Rwpos111_42 in111_42 sp111_42 78000.000000
Rwpos111_43 in111_43 sp111_43 78000.000000
Rwpos111_44 in111_44 sp111_44 202000.000000
Rwpos111_45 in111_45 sp111_45 202000.000000
Rwpos111_46 in111_46 sp111_46 78000.000000
Rwpos111_47 in111_47 sp111_47 202000.000000
Rwpos111_48 in111_48 sp111_48 78000.000000
Rwpos111_49 in111_49 sp111_49 78000.000000
Rwpos111_50 in111_50 sp111_50 78000.000000
Rwpos111_51 in111_51 sp111_51 78000.000000
Rwpos111_52 in111_52 sp111_52 78000.000000
Rwpos111_53 in111_53 sp111_53 202000.000000
Rwpos111_54 in111_54 sp111_54 202000.000000
Rwpos111_55 in111_55 sp111_55 202000.000000
Rwpos111_56 in111_56 sp111_56 78000.000000
Rwpos111_57 in111_57 sp111_57 78000.000000
Rwpos111_58 in111_58 sp111_58 78000.000000
Rwpos111_59 in111_59 sp111_59 78000.000000
Rwpos111_60 in111_60 sp111_60 202000.000000
Rwpos111_61 in111_61 sp111_61 78000.000000
Rwpos111_62 in111_62 sp111_62 78000.000000
Rwpos111_63 in111_63 sp111_63 202000.000000
Rwpos111_64 in111_64 sp111_64 202000.000000
Rwpos111_65 in111_65 sp111_65 78000.000000
Rwpos111_66 in111_66 sp111_66 78000.000000
Rwpos111_67 in111_67 sp111_67 202000.000000
Rwpos111_68 in111_68 sp111_68 202000.000000
Rwpos111_69 in111_69 sp111_69 78000.000000
Rwpos111_70 in111_70 sp111_70 202000.000000
Rwpos111_71 in111_71 sp111_71 202000.000000
Rwpos111_72 in111_72 sp111_72 202000.000000
Rwpos111_73 in111_73 sp111_73 78000.000000
Rwpos111_74 in111_74 sp111_74 78000.000000
Rwpos111_75 in111_75 sp111_75 202000.000000
Rwpos111_76 in111_76 sp111_76 78000.000000
Rwpos111_77 in111_77 sp111_77 202000.000000
Rwpos111_78 in111_78 sp111_78 202000.000000
Rwpos111_79 in111_79 sp111_79 78000.000000
Rwpos111_80 in111_80 sp111_80 202000.000000
Rwpos111_81 in111_81 sp111_81 78000.000000
Rwpos111_82 in111_82 sp111_82 202000.000000
Rwpos111_83 in111_83 sp111_83 202000.000000
Rwpos111_84 in111_84 sp111_84 78000.000000
Rwpos112_1 in112_1 sp112_1 202000.000000
Rwpos112_2 in112_2 sp112_2 78000.000000
Rwpos112_3 in112_3 sp112_3 202000.000000
Rwpos112_4 in112_4 sp112_4 78000.000000
Rwpos112_5 in112_5 sp112_5 202000.000000
Rwpos112_6 in112_6 sp112_6 202000.000000
Rwpos112_7 in112_7 sp112_7 78000.000000
Rwpos112_8 in112_8 sp112_8 202000.000000
Rwpos112_9 in112_9 sp112_9 202000.000000
Rwpos112_10 in112_10 sp112_10 78000.000000
Rwpos112_11 in112_11 sp112_11 202000.000000
Rwpos112_12 in112_12 sp112_12 202000.000000
Rwpos112_13 in112_13 sp112_13 78000.000000
Rwpos112_14 in112_14 sp112_14 78000.000000
Rwpos112_15 in112_15 sp112_15 78000.000000
Rwpos112_16 in112_16 sp112_16 78000.000000
Rwpos112_17 in112_17 sp112_17 202000.000000
Rwpos112_18 in112_18 sp112_18 78000.000000
Rwpos112_19 in112_19 sp112_19 202000.000000
Rwpos112_20 in112_20 sp112_20 78000.000000
Rwpos112_21 in112_21 sp112_21 78000.000000
Rwpos112_22 in112_22 sp112_22 202000.000000
Rwpos112_23 in112_23 sp112_23 78000.000000
Rwpos112_24 in112_24 sp112_24 202000.000000
Rwpos112_25 in112_25 sp112_25 78000.000000
Rwpos112_26 in112_26 sp112_26 78000.000000
Rwpos112_27 in112_27 sp112_27 202000.000000
Rwpos112_28 in112_28 sp112_28 78000.000000
Rwpos112_29 in112_29 sp112_29 78000.000000
Rwpos112_30 in112_30 sp112_30 78000.000000
Rwpos112_31 in112_31 sp112_31 202000.000000
Rwpos112_32 in112_32 sp112_32 202000.000000
Rwpos112_33 in112_33 sp112_33 78000.000000
Rwpos112_34 in112_34 sp112_34 78000.000000
Rwpos112_35 in112_35 sp112_35 202000.000000
Rwpos112_36 in112_36 sp112_36 78000.000000
Rwpos112_37 in112_37 sp112_37 78000.000000
Rwpos112_38 in112_38 sp112_38 202000.000000
Rwpos112_39 in112_39 sp112_39 78000.000000
Rwpos112_40 in112_40 sp112_40 202000.000000
Rwpos112_41 in112_41 sp112_41 78000.000000
Rwpos112_42 in112_42 sp112_42 78000.000000
Rwpos112_43 in112_43 sp112_43 78000.000000
Rwpos112_44 in112_44 sp112_44 78000.000000
Rwpos112_45 in112_45 sp112_45 78000.000000
Rwpos112_46 in112_46 sp112_46 202000.000000
Rwpos112_47 in112_47 sp112_47 78000.000000
Rwpos112_48 in112_48 sp112_48 202000.000000
Rwpos112_49 in112_49 sp112_49 202000.000000
Rwpos112_50 in112_50 sp112_50 78000.000000
Rwpos112_51 in112_51 sp112_51 78000.000000
Rwpos112_52 in112_52 sp112_52 78000.000000
Rwpos112_53 in112_53 sp112_53 202000.000000
Rwpos112_54 in112_54 sp112_54 78000.000000
Rwpos112_55 in112_55 sp112_55 78000.000000
Rwpos112_56 in112_56 sp112_56 78000.000000
Rwpos112_57 in112_57 sp112_57 202000.000000
Rwpos112_58 in112_58 sp112_58 78000.000000
Rwpos112_59 in112_59 sp112_59 202000.000000
Rwpos112_60 in112_60 sp112_60 78000.000000
Rwpos112_61 in112_61 sp112_61 202000.000000
Rwpos112_62 in112_62 sp112_62 78000.000000
Rwpos112_63 in112_63 sp112_63 202000.000000
Rwpos112_64 in112_64 sp112_64 202000.000000
Rwpos112_65 in112_65 sp112_65 78000.000000
Rwpos112_66 in112_66 sp112_66 78000.000000
Rwpos112_67 in112_67 sp112_67 202000.000000
Rwpos112_68 in112_68 sp112_68 78000.000000
Rwpos112_69 in112_69 sp112_69 78000.000000
Rwpos112_70 in112_70 sp112_70 78000.000000
Rwpos112_71 in112_71 sp112_71 78000.000000
Rwpos112_72 in112_72 sp112_72 202000.000000
Rwpos112_73 in112_73 sp112_73 202000.000000
Rwpos112_74 in112_74 sp112_74 202000.000000
Rwpos112_75 in112_75 sp112_75 202000.000000
Rwpos112_76 in112_76 sp112_76 202000.000000
Rwpos112_77 in112_77 sp112_77 78000.000000
Rwpos112_78 in112_78 sp112_78 78000.000000
Rwpos112_79 in112_79 sp112_79 78000.000000
Rwpos112_80 in112_80 sp112_80 78000.000000
Rwpos112_81 in112_81 sp112_81 78000.000000
Rwpos112_82 in112_82 sp112_82 202000.000000
Rwpos112_83 in112_83 sp112_83 78000.000000
Rwpos112_84 in112_84 sp112_84 78000.000000
Rwpos113_1 in113_1 sp113_1 78000.000000
Rwpos113_2 in113_2 sp113_2 202000.000000
Rwpos113_3 in113_3 sp113_3 78000.000000
Rwpos113_4 in113_4 sp113_4 78000.000000
Rwpos113_5 in113_5 sp113_5 78000.000000
Rwpos113_6 in113_6 sp113_6 78000.000000
Rwpos113_7 in113_7 sp113_7 202000.000000
Rwpos113_8 in113_8 sp113_8 78000.000000
Rwpos113_9 in113_9 sp113_9 202000.000000
Rwpos113_10 in113_10 sp113_10 202000.000000
Rwpos113_11 in113_11 sp113_11 78000.000000
Rwpos113_12 in113_12 sp113_12 78000.000000
Rwpos113_13 in113_13 sp113_13 78000.000000
Rwpos113_14 in113_14 sp113_14 78000.000000
Rwpos113_15 in113_15 sp113_15 202000.000000
Rwpos113_16 in113_16 sp113_16 78000.000000
Rwpos113_17 in113_17 sp113_17 78000.000000
Rwpos113_18 in113_18 sp113_18 78000.000000
Rwpos113_19 in113_19 sp113_19 202000.000000
Rwpos113_20 in113_20 sp113_20 78000.000000
Rwpos113_21 in113_21 sp113_21 202000.000000
Rwpos113_22 in113_22 sp113_22 78000.000000
Rwpos113_23 in113_23 sp113_23 78000.000000
Rwpos113_24 in113_24 sp113_24 78000.000000
Rwpos113_25 in113_25 sp113_25 202000.000000
Rwpos113_26 in113_26 sp113_26 202000.000000
Rwpos113_27 in113_27 sp113_27 78000.000000
Rwpos113_28 in113_28 sp113_28 78000.000000
Rwpos113_29 in113_29 sp113_29 202000.000000
Rwpos113_30 in113_30 sp113_30 78000.000000
Rwpos113_31 in113_31 sp113_31 78000.000000
Rwpos113_32 in113_32 sp113_32 202000.000000
Rwpos113_33 in113_33 sp113_33 202000.000000
Rwpos113_34 in113_34 sp113_34 78000.000000
Rwpos113_35 in113_35 sp113_35 78000.000000
Rwpos113_36 in113_36 sp113_36 202000.000000
Rwpos113_37 in113_37 sp113_37 202000.000000
Rwpos113_38 in113_38 sp113_38 202000.000000
Rwpos113_39 in113_39 sp113_39 202000.000000
Rwpos113_40 in113_40 sp113_40 78000.000000
Rwpos113_41 in113_41 sp113_41 78000.000000
Rwpos113_42 in113_42 sp113_42 202000.000000
Rwpos113_43 in113_43 sp113_43 78000.000000
Rwpos113_44 in113_44 sp113_44 78000.000000
Rwpos113_45 in113_45 sp113_45 78000.000000
Rwpos113_46 in113_46 sp113_46 78000.000000
Rwpos113_47 in113_47 sp113_47 202000.000000
Rwpos113_48 in113_48 sp113_48 78000.000000
Rwpos113_49 in113_49 sp113_49 202000.000000
Rwpos113_50 in113_50 sp113_50 202000.000000
Rwpos113_51 in113_51 sp113_51 202000.000000
Rwpos113_52 in113_52 sp113_52 202000.000000
Rwpos113_53 in113_53 sp113_53 202000.000000
Rwpos113_54 in113_54 sp113_54 78000.000000
Rwpos113_55 in113_55 sp113_55 202000.000000
Rwpos113_56 in113_56 sp113_56 78000.000000
Rwpos113_57 in113_57 sp113_57 78000.000000
Rwpos113_58 in113_58 sp113_58 78000.000000
Rwpos113_59 in113_59 sp113_59 78000.000000
Rwpos113_60 in113_60 sp113_60 202000.000000
Rwpos113_61 in113_61 sp113_61 202000.000000
Rwpos113_62 in113_62 sp113_62 78000.000000
Rwpos113_63 in113_63 sp113_63 202000.000000
Rwpos113_64 in113_64 sp113_64 78000.000000
Rwpos113_65 in113_65 sp113_65 78000.000000
Rwpos113_66 in113_66 sp113_66 202000.000000
Rwpos113_67 in113_67 sp113_67 202000.000000
Rwpos113_68 in113_68 sp113_68 78000.000000
Rwpos113_69 in113_69 sp113_69 78000.000000
Rwpos113_70 in113_70 sp113_70 78000.000000
Rwpos113_71 in113_71 sp113_71 78000.000000
Rwpos113_72 in113_72 sp113_72 78000.000000
Rwpos113_73 in113_73 sp113_73 78000.000000
Rwpos113_74 in113_74 sp113_74 202000.000000
Rwpos113_75 in113_75 sp113_75 78000.000000
Rwpos113_76 in113_76 sp113_76 202000.000000
Rwpos113_77 in113_77 sp113_77 78000.000000
Rwpos113_78 in113_78 sp113_78 202000.000000
Rwpos113_79 in113_79 sp113_79 202000.000000
Rwpos113_80 in113_80 sp113_80 78000.000000
Rwpos113_81 in113_81 sp113_81 78000.000000
Rwpos113_82 in113_82 sp113_82 202000.000000
Rwpos113_83 in113_83 sp113_83 202000.000000
Rwpos113_84 in113_84 sp113_84 202000.000000
Rwpos114_1 in114_1 sp114_1 202000.000000
Rwpos114_2 in114_2 sp114_2 78000.000000
Rwpos114_3 in114_3 sp114_3 78000.000000
Rwpos114_4 in114_4 sp114_4 78000.000000
Rwpos114_5 in114_5 sp114_5 202000.000000
Rwpos114_6 in114_6 sp114_6 78000.000000
Rwpos114_7 in114_7 sp114_7 78000.000000
Rwpos114_8 in114_8 sp114_8 202000.000000
Rwpos114_9 in114_9 sp114_9 202000.000000
Rwpos114_10 in114_10 sp114_10 78000.000000
Rwpos114_11 in114_11 sp114_11 78000.000000
Rwpos114_12 in114_12 sp114_12 202000.000000
Rwpos114_13 in114_13 sp114_13 78000.000000
Rwpos114_14 in114_14 sp114_14 78000.000000
Rwpos114_15 in114_15 sp114_15 78000.000000
Rwpos114_16 in114_16 sp114_16 78000.000000
Rwpos114_17 in114_17 sp114_17 202000.000000
Rwpos114_18 in114_18 sp114_18 202000.000000
Rwpos114_19 in114_19 sp114_19 78000.000000
Rwpos114_20 in114_20 sp114_20 78000.000000
Rwpos114_21 in114_21 sp114_21 78000.000000
Rwpos114_22 in114_22 sp114_22 78000.000000
Rwpos114_23 in114_23 sp114_23 78000.000000
Rwpos114_24 in114_24 sp114_24 202000.000000
Rwpos114_25 in114_25 sp114_25 78000.000000
Rwpos114_26 in114_26 sp114_26 78000.000000
Rwpos114_27 in114_27 sp114_27 202000.000000
Rwpos114_28 in114_28 sp114_28 78000.000000
Rwpos114_29 in114_29 sp114_29 78000.000000
Rwpos114_30 in114_30 sp114_30 78000.000000
Rwpos114_31 in114_31 sp114_31 78000.000000
Rwpos114_32 in114_32 sp114_32 202000.000000
Rwpos114_33 in114_33 sp114_33 78000.000000
Rwpos114_34 in114_34 sp114_34 202000.000000
Rwpos114_35 in114_35 sp114_35 78000.000000
Rwpos114_36 in114_36 sp114_36 202000.000000
Rwpos114_37 in114_37 sp114_37 78000.000000
Rwpos114_38 in114_38 sp114_38 78000.000000
Rwpos114_39 in114_39 sp114_39 202000.000000
Rwpos114_40 in114_40 sp114_40 78000.000000
Rwpos114_41 in114_41 sp114_41 202000.000000
Rwpos114_42 in114_42 sp114_42 78000.000000
Rwpos114_43 in114_43 sp114_43 78000.000000
Rwpos114_44 in114_44 sp114_44 202000.000000
Rwpos114_45 in114_45 sp114_45 78000.000000
Rwpos114_46 in114_46 sp114_46 78000.000000
Rwpos114_47 in114_47 sp114_47 78000.000000
Rwpos114_48 in114_48 sp114_48 78000.000000
Rwpos114_49 in114_49 sp114_49 78000.000000
Rwpos114_50 in114_50 sp114_50 78000.000000
Rwpos114_51 in114_51 sp114_51 78000.000000
Rwpos114_52 in114_52 sp114_52 78000.000000
Rwpos114_53 in114_53 sp114_53 78000.000000
Rwpos114_54 in114_54 sp114_54 78000.000000
Rwpos114_55 in114_55 sp114_55 78000.000000
Rwpos114_56 in114_56 sp114_56 202000.000000
Rwpos114_57 in114_57 sp114_57 202000.000000
Rwpos114_58 in114_58 sp114_58 78000.000000
Rwpos114_59 in114_59 sp114_59 78000.000000
Rwpos114_60 in114_60 sp114_60 202000.000000
Rwpos114_61 in114_61 sp114_61 202000.000000
Rwpos114_62 in114_62 sp114_62 78000.000000
Rwpos114_63 in114_63 sp114_63 78000.000000
Rwpos114_64 in114_64 sp114_64 202000.000000
Rwpos114_65 in114_65 sp114_65 78000.000000
Rwpos114_66 in114_66 sp114_66 78000.000000
Rwpos114_67 in114_67 sp114_67 78000.000000
Rwpos114_68 in114_68 sp114_68 202000.000000
Rwpos114_69 in114_69 sp114_69 202000.000000
Rwpos114_70 in114_70 sp114_70 78000.000000
Rwpos114_71 in114_71 sp114_71 202000.000000
Rwpos114_72 in114_72 sp114_72 78000.000000
Rwpos114_73 in114_73 sp114_73 202000.000000
Rwpos114_74 in114_74 sp114_74 202000.000000
Rwpos114_75 in114_75 sp114_75 202000.000000
Rwpos114_76 in114_76 sp114_76 78000.000000
Rwpos114_77 in114_77 sp114_77 202000.000000
Rwpos114_78 in114_78 sp114_78 202000.000000
Rwpos114_79 in114_79 sp114_79 202000.000000
Rwpos114_80 in114_80 sp114_80 202000.000000
Rwpos114_81 in114_81 sp114_81 78000.000000
Rwpos114_82 in114_82 sp114_82 202000.000000
Rwpos114_83 in114_83 sp114_83 202000.000000
Rwpos114_84 in114_84 sp114_84 78000.000000
Rwpos115_1 in115_1 sp115_1 78000.000000
Rwpos115_2 in115_2 sp115_2 78000.000000
Rwpos115_3 in115_3 sp115_3 78000.000000
Rwpos115_4 in115_4 sp115_4 202000.000000
Rwpos115_5 in115_5 sp115_5 78000.000000
Rwpos115_6 in115_6 sp115_6 78000.000000
Rwpos115_7 in115_7 sp115_7 202000.000000
Rwpos115_8 in115_8 sp115_8 78000.000000
Rwpos115_9 in115_9 sp115_9 78000.000000
Rwpos115_10 in115_10 sp115_10 202000.000000
Rwpos115_11 in115_11 sp115_11 78000.000000
Rwpos115_12 in115_12 sp115_12 202000.000000
Rwpos115_13 in115_13 sp115_13 202000.000000
Rwpos115_14 in115_14 sp115_14 202000.000000
Rwpos115_15 in115_15 sp115_15 78000.000000
Rwpos115_16 in115_16 sp115_16 202000.000000
Rwpos115_17 in115_17 sp115_17 78000.000000
Rwpos115_18 in115_18 sp115_18 202000.000000
Rwpos115_19 in115_19 sp115_19 78000.000000
Rwpos115_20 in115_20 sp115_20 202000.000000
Rwpos115_21 in115_21 sp115_21 78000.000000
Rwpos115_22 in115_22 sp115_22 78000.000000
Rwpos115_23 in115_23 sp115_23 202000.000000
Rwpos115_24 in115_24 sp115_24 78000.000000
Rwpos115_25 in115_25 sp115_25 78000.000000
Rwpos115_26 in115_26 sp115_26 202000.000000
Rwpos115_27 in115_27 sp115_27 78000.000000
Rwpos115_28 in115_28 sp115_28 202000.000000
Rwpos115_29 in115_29 sp115_29 78000.000000
Rwpos115_30 in115_30 sp115_30 78000.000000
Rwpos115_31 in115_31 sp115_31 78000.000000
Rwpos115_32 in115_32 sp115_32 202000.000000
Rwpos115_33 in115_33 sp115_33 78000.000000
Rwpos115_34 in115_34 sp115_34 202000.000000
Rwpos115_35 in115_35 sp115_35 202000.000000
Rwpos115_36 in115_36 sp115_36 78000.000000
Rwpos115_37 in115_37 sp115_37 202000.000000
Rwpos115_38 in115_38 sp115_38 202000.000000
Rwpos115_39 in115_39 sp115_39 202000.000000
Rwpos115_40 in115_40 sp115_40 202000.000000
Rwpos115_41 in115_41 sp115_41 202000.000000
Rwpos115_42 in115_42 sp115_42 202000.000000
Rwpos115_43 in115_43 sp115_43 78000.000000
Rwpos115_44 in115_44 sp115_44 78000.000000
Rwpos115_45 in115_45 sp115_45 202000.000000
Rwpos115_46 in115_46 sp115_46 78000.000000
Rwpos115_47 in115_47 sp115_47 202000.000000
Rwpos115_48 in115_48 sp115_48 202000.000000
Rwpos115_49 in115_49 sp115_49 202000.000000
Rwpos115_50 in115_50 sp115_50 202000.000000
Rwpos115_51 in115_51 sp115_51 202000.000000
Rwpos115_52 in115_52 sp115_52 202000.000000
Rwpos115_53 in115_53 sp115_53 78000.000000
Rwpos115_54 in115_54 sp115_54 78000.000000
Rwpos115_55 in115_55 sp115_55 202000.000000
Rwpos115_56 in115_56 sp115_56 78000.000000
Rwpos115_57 in115_57 sp115_57 78000.000000
Rwpos115_58 in115_58 sp115_58 78000.000000
Rwpos115_59 in115_59 sp115_59 78000.000000
Rwpos115_60 in115_60 sp115_60 78000.000000
Rwpos115_61 in115_61 sp115_61 78000.000000
Rwpos115_62 in115_62 sp115_62 202000.000000
Rwpos115_63 in115_63 sp115_63 202000.000000
Rwpos115_64 in115_64 sp115_64 78000.000000
Rwpos115_65 in115_65 sp115_65 78000.000000
Rwpos115_66 in115_66 sp115_66 78000.000000
Rwpos115_67 in115_67 sp115_67 78000.000000
Rwpos115_68 in115_68 sp115_68 202000.000000
Rwpos115_69 in115_69 sp115_69 202000.000000
Rwpos115_70 in115_70 sp115_70 202000.000000
Rwpos115_71 in115_71 sp115_71 202000.000000
Rwpos115_72 in115_72 sp115_72 202000.000000
Rwpos115_73 in115_73 sp115_73 78000.000000
Rwpos115_74 in115_74 sp115_74 78000.000000
Rwpos115_75 in115_75 sp115_75 202000.000000
Rwpos115_76 in115_76 sp115_76 78000.000000
Rwpos115_77 in115_77 sp115_77 202000.000000
Rwpos115_78 in115_78 sp115_78 78000.000000
Rwpos115_79 in115_79 sp115_79 202000.000000
Rwpos115_80 in115_80 sp115_80 202000.000000
Rwpos115_81 in115_81 sp115_81 202000.000000
Rwpos115_82 in115_82 sp115_82 78000.000000
Rwpos115_83 in115_83 sp115_83 78000.000000
Rwpos115_84 in115_84 sp115_84 202000.000000
Rwpos116_1 in116_1 sp116_1 78000.000000
Rwpos116_2 in116_2 sp116_2 202000.000000
Rwpos116_3 in116_3 sp116_3 202000.000000
Rwpos116_4 in116_4 sp116_4 78000.000000
Rwpos116_5 in116_5 sp116_5 78000.000000
Rwpos116_6 in116_6 sp116_6 202000.000000
Rwpos116_7 in116_7 sp116_7 202000.000000
Rwpos116_8 in116_8 sp116_8 202000.000000
Rwpos116_9 in116_9 sp116_9 78000.000000
Rwpos116_10 in116_10 sp116_10 202000.000000
Rwpos116_11 in116_11 sp116_11 78000.000000
Rwpos116_12 in116_12 sp116_12 78000.000000
Rwpos116_13 in116_13 sp116_13 202000.000000
Rwpos116_14 in116_14 sp116_14 78000.000000
Rwpos116_15 in116_15 sp116_15 78000.000000
Rwpos116_16 in116_16 sp116_16 202000.000000
Rwpos116_17 in116_17 sp116_17 202000.000000
Rwpos116_18 in116_18 sp116_18 78000.000000
Rwpos116_19 in116_19 sp116_19 202000.000000
Rwpos116_20 in116_20 sp116_20 202000.000000
Rwpos116_21 in116_21 sp116_21 202000.000000
Rwpos116_22 in116_22 sp116_22 202000.000000
Rwpos116_23 in116_23 sp116_23 78000.000000
Rwpos116_24 in116_24 sp116_24 202000.000000
Rwpos116_25 in116_25 sp116_25 202000.000000
Rwpos116_26 in116_26 sp116_26 202000.000000
Rwpos116_27 in116_27 sp116_27 202000.000000
Rwpos116_28 in116_28 sp116_28 78000.000000
Rwpos116_29 in116_29 sp116_29 78000.000000
Rwpos116_30 in116_30 sp116_30 202000.000000
Rwpos116_31 in116_31 sp116_31 78000.000000
Rwpos116_32 in116_32 sp116_32 78000.000000
Rwpos116_33 in116_33 sp116_33 202000.000000
Rwpos116_34 in116_34 sp116_34 78000.000000
Rwpos116_35 in116_35 sp116_35 78000.000000
Rwpos116_36 in116_36 sp116_36 78000.000000
Rwpos116_37 in116_37 sp116_37 78000.000000
Rwpos116_38 in116_38 sp116_38 202000.000000
Rwpos116_39 in116_39 sp116_39 78000.000000
Rwpos116_40 in116_40 sp116_40 78000.000000
Rwpos116_41 in116_41 sp116_41 202000.000000
Rwpos116_42 in116_42 sp116_42 202000.000000
Rwpos116_43 in116_43 sp116_43 78000.000000
Rwpos116_44 in116_44 sp116_44 202000.000000
Rwpos116_45 in116_45 sp116_45 202000.000000
Rwpos116_46 in116_46 sp116_46 78000.000000
Rwpos116_47 in116_47 sp116_47 78000.000000
Rwpos116_48 in116_48 sp116_48 202000.000000
Rwpos116_49 in116_49 sp116_49 78000.000000
Rwpos116_50 in116_50 sp116_50 78000.000000
Rwpos116_51 in116_51 sp116_51 78000.000000
Rwpos116_52 in116_52 sp116_52 78000.000000
Rwpos116_53 in116_53 sp116_53 78000.000000
Rwpos116_54 in116_54 sp116_54 202000.000000
Rwpos116_55 in116_55 sp116_55 78000.000000
Rwpos116_56 in116_56 sp116_56 78000.000000
Rwpos116_57 in116_57 sp116_57 78000.000000
Rwpos116_58 in116_58 sp116_58 78000.000000
Rwpos116_59 in116_59 sp116_59 78000.000000
Rwpos116_60 in116_60 sp116_60 202000.000000
Rwpos116_61 in116_61 sp116_61 78000.000000
Rwpos116_62 in116_62 sp116_62 78000.000000
Rwpos116_63 in116_63 sp116_63 202000.000000
Rwpos116_64 in116_64 sp116_64 202000.000000
Rwpos116_65 in116_65 sp116_65 202000.000000
Rwpos116_66 in116_66 sp116_66 78000.000000
Rwpos116_67 in116_67 sp116_67 78000.000000
Rwpos116_68 in116_68 sp116_68 78000.000000
Rwpos116_69 in116_69 sp116_69 78000.000000
Rwpos116_70 in116_70 sp116_70 202000.000000
Rwpos116_71 in116_71 sp116_71 78000.000000
Rwpos116_72 in116_72 sp116_72 202000.000000
Rwpos116_73 in116_73 sp116_73 78000.000000
Rwpos116_74 in116_74 sp116_74 202000.000000
Rwpos116_75 in116_75 sp116_75 78000.000000
Rwpos116_76 in116_76 sp116_76 78000.000000
Rwpos116_77 in116_77 sp116_77 78000.000000
Rwpos116_78 in116_78 sp116_78 78000.000000
Rwpos116_79 in116_79 sp116_79 78000.000000
Rwpos116_80 in116_80 sp116_80 78000.000000
Rwpos116_81 in116_81 sp116_81 202000.000000
Rwpos116_82 in116_82 sp116_82 78000.000000
Rwpos116_83 in116_83 sp116_83 202000.000000
Rwpos116_84 in116_84 sp116_84 202000.000000
Rwpos117_1 in117_1 sp117_1 78000.000000
Rwpos117_2 in117_2 sp117_2 78000.000000
Rwpos117_3 in117_3 sp117_3 202000.000000
Rwpos117_4 in117_4 sp117_4 202000.000000
Rwpos117_5 in117_5 sp117_5 78000.000000
Rwpos117_6 in117_6 sp117_6 202000.000000
Rwpos117_7 in117_7 sp117_7 78000.000000
Rwpos117_8 in117_8 sp117_8 78000.000000
Rwpos117_9 in117_9 sp117_9 78000.000000
Rwpos117_10 in117_10 sp117_10 78000.000000
Rwpos117_11 in117_11 sp117_11 202000.000000
Rwpos117_12 in117_12 sp117_12 78000.000000
Rwpos117_13 in117_13 sp117_13 78000.000000
Rwpos117_14 in117_14 sp117_14 202000.000000
Rwpos117_15 in117_15 sp117_15 202000.000000
Rwpos117_16 in117_16 sp117_16 78000.000000
Rwpos117_17 in117_17 sp117_17 202000.000000
Rwpos117_18 in117_18 sp117_18 202000.000000
Rwpos117_19 in117_19 sp117_19 202000.000000
Rwpos117_20 in117_20 sp117_20 78000.000000
Rwpos117_21 in117_21 sp117_21 78000.000000
Rwpos117_22 in117_22 sp117_22 202000.000000
Rwpos117_23 in117_23 sp117_23 202000.000000
Rwpos117_24 in117_24 sp117_24 202000.000000
Rwpos117_25 in117_25 sp117_25 78000.000000
Rwpos117_26 in117_26 sp117_26 78000.000000
Rwpos117_27 in117_27 sp117_27 78000.000000
Rwpos117_28 in117_28 sp117_28 78000.000000
Rwpos117_29 in117_29 sp117_29 202000.000000
Rwpos117_30 in117_30 sp117_30 78000.000000
Rwpos117_31 in117_31 sp117_31 202000.000000
Rwpos117_32 in117_32 sp117_32 78000.000000
Rwpos117_33 in117_33 sp117_33 78000.000000
Rwpos117_34 in117_34 sp117_34 202000.000000
Rwpos117_35 in117_35 sp117_35 78000.000000
Rwpos117_36 in117_36 sp117_36 202000.000000
Rwpos117_37 in117_37 sp117_37 78000.000000
Rwpos117_38 in117_38 sp117_38 202000.000000
Rwpos117_39 in117_39 sp117_39 202000.000000
Rwpos117_40 in117_40 sp117_40 202000.000000
Rwpos117_41 in117_41 sp117_41 202000.000000
Rwpos117_42 in117_42 sp117_42 78000.000000
Rwpos117_43 in117_43 sp117_43 78000.000000
Rwpos117_44 in117_44 sp117_44 78000.000000
Rwpos117_45 in117_45 sp117_45 78000.000000
Rwpos117_46 in117_46 sp117_46 202000.000000
Rwpos117_47 in117_47 sp117_47 78000.000000
Rwpos117_48 in117_48 sp117_48 202000.000000
Rwpos117_49 in117_49 sp117_49 202000.000000
Rwpos117_50 in117_50 sp117_50 78000.000000
Rwpos117_51 in117_51 sp117_51 78000.000000
Rwpos117_52 in117_52 sp117_52 78000.000000
Rwpos117_53 in117_53 sp117_53 202000.000000
Rwpos117_54 in117_54 sp117_54 78000.000000
Rwpos117_55 in117_55 sp117_55 78000.000000
Rwpos117_56 in117_56 sp117_56 202000.000000
Rwpos117_57 in117_57 sp117_57 202000.000000
Rwpos117_58 in117_58 sp117_58 202000.000000
Rwpos117_59 in117_59 sp117_59 78000.000000
Rwpos117_60 in117_60 sp117_60 78000.000000
Rwpos117_61 in117_61 sp117_61 78000.000000
Rwpos117_62 in117_62 sp117_62 78000.000000
Rwpos117_63 in117_63 sp117_63 78000.000000
Rwpos117_64 in117_64 sp117_64 78000.000000
Rwpos117_65 in117_65 sp117_65 202000.000000
Rwpos117_66 in117_66 sp117_66 78000.000000
Rwpos117_67 in117_67 sp117_67 202000.000000
Rwpos117_68 in117_68 sp117_68 202000.000000
Rwpos117_69 in117_69 sp117_69 78000.000000
Rwpos117_70 in117_70 sp117_70 202000.000000
Rwpos117_71 in117_71 sp117_71 202000.000000
Rwpos117_72 in117_72 sp117_72 78000.000000
Rwpos117_73 in117_73 sp117_73 78000.000000
Rwpos117_74 in117_74 sp117_74 78000.000000
Rwpos117_75 in117_75 sp117_75 202000.000000
Rwpos117_76 in117_76 sp117_76 78000.000000
Rwpos117_77 in117_77 sp117_77 202000.000000
Rwpos117_78 in117_78 sp117_78 202000.000000
Rwpos117_79 in117_79 sp117_79 202000.000000
Rwpos117_80 in117_80 sp117_80 78000.000000
Rwpos117_81 in117_81 sp117_81 78000.000000
Rwpos117_82 in117_82 sp117_82 78000.000000
Rwpos117_83 in117_83 sp117_83 78000.000000
Rwpos117_84 in117_84 sp117_84 202000.000000
Rwpos118_1 in118_1 sp118_1 202000.000000
Rwpos118_2 in118_2 sp118_2 202000.000000
Rwpos118_3 in118_3 sp118_3 78000.000000
Rwpos118_4 in118_4 sp118_4 78000.000000
Rwpos118_5 in118_5 sp118_5 78000.000000
Rwpos118_6 in118_6 sp118_6 78000.000000
Rwpos118_7 in118_7 sp118_7 202000.000000
Rwpos118_8 in118_8 sp118_8 202000.000000
Rwpos118_9 in118_9 sp118_9 202000.000000
Rwpos118_10 in118_10 sp118_10 78000.000000
Rwpos118_11 in118_11 sp118_11 78000.000000
Rwpos118_12 in118_12 sp118_12 78000.000000
Rwpos118_13 in118_13 sp118_13 78000.000000
Rwpos118_14 in118_14 sp118_14 78000.000000
Rwpos118_15 in118_15 sp118_15 202000.000000
Rwpos118_16 in118_16 sp118_16 78000.000000
Rwpos118_17 in118_17 sp118_17 78000.000000
Rwpos118_18 in118_18 sp118_18 78000.000000
Rwpos118_19 in118_19 sp118_19 78000.000000
Rwpos118_20 in118_20 sp118_20 78000.000000
Rwpos118_21 in118_21 sp118_21 78000.000000
Rwpos118_22 in118_22 sp118_22 202000.000000
Rwpos118_23 in118_23 sp118_23 78000.000000
Rwpos118_24 in118_24 sp118_24 202000.000000
Rwpos118_25 in118_25 sp118_25 202000.000000
Rwpos118_26 in118_26 sp118_26 202000.000000
Rwpos118_27 in118_27 sp118_27 202000.000000
Rwpos118_28 in118_28 sp118_28 202000.000000
Rwpos118_29 in118_29 sp118_29 78000.000000
Rwpos118_30 in118_30 sp118_30 202000.000000
Rwpos118_31 in118_31 sp118_31 78000.000000
Rwpos118_32 in118_32 sp118_32 78000.000000
Rwpos118_33 in118_33 sp118_33 78000.000000
Rwpos118_34 in118_34 sp118_34 78000.000000
Rwpos118_35 in118_35 sp118_35 202000.000000
Rwpos118_36 in118_36 sp118_36 202000.000000
Rwpos118_37 in118_37 sp118_37 78000.000000
Rwpos118_38 in118_38 sp118_38 78000.000000
Rwpos118_39 in118_39 sp118_39 202000.000000
Rwpos118_40 in118_40 sp118_40 78000.000000
Rwpos118_41 in118_41 sp118_41 202000.000000
Rwpos118_42 in118_42 sp118_42 202000.000000
Rwpos118_43 in118_43 sp118_43 78000.000000
Rwpos118_44 in118_44 sp118_44 202000.000000
Rwpos118_45 in118_45 sp118_45 78000.000000
Rwpos118_46 in118_46 sp118_46 78000.000000
Rwpos118_47 in118_47 sp118_47 202000.000000
Rwpos118_48 in118_48 sp118_48 78000.000000
Rwpos118_49 in118_49 sp118_49 202000.000000
Rwpos118_50 in118_50 sp118_50 78000.000000
Rwpos118_51 in118_51 sp118_51 78000.000000
Rwpos118_52 in118_52 sp118_52 202000.000000
Rwpos118_53 in118_53 sp118_53 78000.000000
Rwpos118_54 in118_54 sp118_54 202000.000000
Rwpos118_55 in118_55 sp118_55 202000.000000
Rwpos118_56 in118_56 sp118_56 78000.000000
Rwpos118_57 in118_57 sp118_57 202000.000000
Rwpos118_58 in118_58 sp118_58 78000.000000
Rwpos118_59 in118_59 sp118_59 78000.000000
Rwpos118_60 in118_60 sp118_60 202000.000000
Rwpos118_61 in118_61 sp118_61 78000.000000
Rwpos118_62 in118_62 sp118_62 78000.000000
Rwpos118_63 in118_63 sp118_63 202000.000000
Rwpos118_64 in118_64 sp118_64 78000.000000
Rwpos118_65 in118_65 sp118_65 202000.000000
Rwpos118_66 in118_66 sp118_66 78000.000000
Rwpos118_67 in118_67 sp118_67 78000.000000
Rwpos118_68 in118_68 sp118_68 78000.000000
Rwpos118_69 in118_69 sp118_69 78000.000000
Rwpos118_70 in118_70 sp118_70 202000.000000
Rwpos118_71 in118_71 sp118_71 78000.000000
Rwpos118_72 in118_72 sp118_72 202000.000000
Rwpos118_73 in118_73 sp118_73 78000.000000
Rwpos118_74 in118_74 sp118_74 202000.000000
Rwpos118_75 in118_75 sp118_75 78000.000000
Rwpos118_76 in118_76 sp118_76 202000.000000
Rwpos118_77 in118_77 sp118_77 78000.000000
Rwpos118_78 in118_78 sp118_78 202000.000000
Rwpos118_79 in118_79 sp118_79 78000.000000
Rwpos118_80 in118_80 sp118_80 78000.000000
Rwpos118_81 in118_81 sp118_81 78000.000000
Rwpos118_82 in118_82 sp118_82 202000.000000
Rwpos118_83 in118_83 sp118_83 78000.000000
Rwpos118_84 in118_84 sp118_84 78000.000000
Rwpos119_1 in119_1 sp119_1 202000.000000
Rwpos119_2 in119_2 sp119_2 78000.000000
Rwpos119_3 in119_3 sp119_3 202000.000000
Rwpos119_4 in119_4 sp119_4 202000.000000
Rwpos119_5 in119_5 sp119_5 202000.000000
Rwpos119_6 in119_6 sp119_6 202000.000000
Rwpos119_7 in119_7 sp119_7 78000.000000
Rwpos119_8 in119_8 sp119_8 202000.000000
Rwpos119_9 in119_9 sp119_9 78000.000000
Rwpos119_10 in119_10 sp119_10 202000.000000
Rwpos119_11 in119_11 sp119_11 78000.000000
Rwpos119_12 in119_12 sp119_12 202000.000000
Rwpos119_13 in119_13 sp119_13 202000.000000
Rwpos119_14 in119_14 sp119_14 202000.000000
Rwpos119_15 in119_15 sp119_15 78000.000000
Rwpos119_16 in119_16 sp119_16 78000.000000
Rwpos119_17 in119_17 sp119_17 78000.000000
Rwpos119_18 in119_18 sp119_18 202000.000000
Rwpos119_19 in119_19 sp119_19 78000.000000
Rwpos119_20 in119_20 sp119_20 202000.000000
Rwpos119_21 in119_21 sp119_21 78000.000000
Rwpos119_22 in119_22 sp119_22 78000.000000
Rwpos119_23 in119_23 sp119_23 78000.000000
Rwpos119_24 in119_24 sp119_24 78000.000000
Rwpos119_25 in119_25 sp119_25 78000.000000
Rwpos119_26 in119_26 sp119_26 202000.000000
Rwpos119_27 in119_27 sp119_27 202000.000000
Rwpos119_28 in119_28 sp119_28 202000.000000
Rwpos119_29 in119_29 sp119_29 78000.000000
Rwpos119_30 in119_30 sp119_30 78000.000000
Rwpos119_31 in119_31 sp119_31 202000.000000
Rwpos119_32 in119_32 sp119_32 78000.000000
Rwpos119_33 in119_33 sp119_33 202000.000000
Rwpos119_34 in119_34 sp119_34 78000.000000
Rwpos119_35 in119_35 sp119_35 202000.000000
Rwpos119_36 in119_36 sp119_36 78000.000000
Rwpos119_37 in119_37 sp119_37 78000.000000
Rwpos119_38 in119_38 sp119_38 78000.000000
Rwpos119_39 in119_39 sp119_39 202000.000000
Rwpos119_40 in119_40 sp119_40 78000.000000
Rwpos119_41 in119_41 sp119_41 78000.000000
Rwpos119_42 in119_42 sp119_42 202000.000000
Rwpos119_43 in119_43 sp119_43 78000.000000
Rwpos119_44 in119_44 sp119_44 78000.000000
Rwpos119_45 in119_45 sp119_45 78000.000000
Rwpos119_46 in119_46 sp119_46 202000.000000
Rwpos119_47 in119_47 sp119_47 202000.000000
Rwpos119_48 in119_48 sp119_48 78000.000000
Rwpos119_49 in119_49 sp119_49 78000.000000
Rwpos119_50 in119_50 sp119_50 78000.000000
Rwpos119_51 in119_51 sp119_51 202000.000000
Rwpos119_52 in119_52 sp119_52 78000.000000
Rwpos119_53 in119_53 sp119_53 202000.000000
Rwpos119_54 in119_54 sp119_54 202000.000000
Rwpos119_55 in119_55 sp119_55 202000.000000
Rwpos119_56 in119_56 sp119_56 78000.000000
Rwpos119_57 in119_57 sp119_57 78000.000000
Rwpos119_58 in119_58 sp119_58 78000.000000
Rwpos119_59 in119_59 sp119_59 202000.000000
Rwpos119_60 in119_60 sp119_60 78000.000000
Rwpos119_61 in119_61 sp119_61 78000.000000
Rwpos119_62 in119_62 sp119_62 202000.000000
Rwpos119_63 in119_63 sp119_63 202000.000000
Rwpos119_64 in119_64 sp119_64 78000.000000
Rwpos119_65 in119_65 sp119_65 78000.000000
Rwpos119_66 in119_66 sp119_66 202000.000000
Rwpos119_67 in119_67 sp119_67 202000.000000
Rwpos119_68 in119_68 sp119_68 78000.000000
Rwpos119_69 in119_69 sp119_69 202000.000000
Rwpos119_70 in119_70 sp119_70 202000.000000
Rwpos119_71 in119_71 sp119_71 202000.000000
Rwpos119_72 in119_72 sp119_72 78000.000000
Rwpos119_73 in119_73 sp119_73 78000.000000
Rwpos119_74 in119_74 sp119_74 78000.000000
Rwpos119_75 in119_75 sp119_75 202000.000000
Rwpos119_76 in119_76 sp119_76 202000.000000
Rwpos119_77 in119_77 sp119_77 78000.000000
Rwpos119_78 in119_78 sp119_78 78000.000000
Rwpos119_79 in119_79 sp119_79 78000.000000
Rwpos119_80 in119_80 sp119_80 202000.000000
Rwpos119_81 in119_81 sp119_81 202000.000000
Rwpos119_82 in119_82 sp119_82 78000.000000
Rwpos119_83 in119_83 sp119_83 78000.000000
Rwpos119_84 in119_84 sp119_84 202000.000000
Rwpos120_1 in120_1 sp120_1 78000.000000
Rwpos120_2 in120_2 sp120_2 202000.000000
Rwpos120_3 in120_3 sp120_3 78000.000000
Rwpos120_4 in120_4 sp120_4 78000.000000
Rwpos120_5 in120_5 sp120_5 78000.000000
Rwpos120_6 in120_6 sp120_6 202000.000000
Rwpos120_7 in120_7 sp120_7 202000.000000
Rwpos120_8 in120_8 sp120_8 202000.000000
Rwpos120_9 in120_9 sp120_9 202000.000000
Rwpos120_10 in120_10 sp120_10 202000.000000
Rwpos120_11 in120_11 sp120_11 78000.000000
Rwpos120_12 in120_12 sp120_12 202000.000000
Rwpos120_13 in120_13 sp120_13 78000.000000
Rwpos120_14 in120_14 sp120_14 78000.000000
Rwpos120_15 in120_15 sp120_15 202000.000000
Rwpos120_16 in120_16 sp120_16 78000.000000
Rwpos120_17 in120_17 sp120_17 78000.000000
Rwpos120_18 in120_18 sp120_18 202000.000000
Rwpos120_19 in120_19 sp120_19 78000.000000
Rwpos120_20 in120_20 sp120_20 202000.000000
Rwpos120_21 in120_21 sp120_21 78000.000000
Rwpos120_22 in120_22 sp120_22 78000.000000
Rwpos120_23 in120_23 sp120_23 202000.000000
Rwpos120_24 in120_24 sp120_24 202000.000000
Rwpos120_25 in120_25 sp120_25 78000.000000
Rwpos120_26 in120_26 sp120_26 202000.000000
Rwpos120_27 in120_27 sp120_27 78000.000000
Rwpos120_28 in120_28 sp120_28 78000.000000
Rwpos120_29 in120_29 sp120_29 202000.000000
Rwpos120_30 in120_30 sp120_30 78000.000000
Rwpos120_31 in120_31 sp120_31 78000.000000
Rwpos120_32 in120_32 sp120_32 78000.000000
Rwpos120_33 in120_33 sp120_33 78000.000000
Rwpos120_34 in120_34 sp120_34 202000.000000
Rwpos120_35 in120_35 sp120_35 78000.000000
Rwpos120_36 in120_36 sp120_36 202000.000000
Rwpos120_37 in120_37 sp120_37 202000.000000
Rwpos120_38 in120_38 sp120_38 78000.000000
Rwpos120_39 in120_39 sp120_39 202000.000000
Rwpos120_40 in120_40 sp120_40 202000.000000
Rwpos120_41 in120_41 sp120_41 202000.000000
Rwpos120_42 in120_42 sp120_42 202000.000000
Rwpos120_43 in120_43 sp120_43 78000.000000
Rwpos120_44 in120_44 sp120_44 78000.000000
Rwpos120_45 in120_45 sp120_45 202000.000000
Rwpos120_46 in120_46 sp120_46 202000.000000
Rwpos120_47 in120_47 sp120_47 202000.000000
Rwpos120_48 in120_48 sp120_48 202000.000000
Rwpos120_49 in120_49 sp120_49 202000.000000
Rwpos120_50 in120_50 sp120_50 202000.000000
Rwpos120_51 in120_51 sp120_51 202000.000000
Rwpos120_52 in120_52 sp120_52 202000.000000
Rwpos120_53 in120_53 sp120_53 202000.000000
Rwpos120_54 in120_54 sp120_54 78000.000000
Rwpos120_55 in120_55 sp120_55 202000.000000
Rwpos120_56 in120_56 sp120_56 78000.000000
Rwpos120_57 in120_57 sp120_57 78000.000000
Rwpos120_58 in120_58 sp120_58 78000.000000
Rwpos120_59 in120_59 sp120_59 78000.000000
Rwpos120_60 in120_60 sp120_60 202000.000000
Rwpos120_61 in120_61 sp120_61 78000.000000
Rwpos120_62 in120_62 sp120_62 202000.000000
Rwpos120_63 in120_63 sp120_63 202000.000000
Rwpos120_64 in120_64 sp120_64 202000.000000
Rwpos120_65 in120_65 sp120_65 78000.000000
Rwpos120_66 in120_66 sp120_66 202000.000000
Rwpos120_67 in120_67 sp120_67 202000.000000
Rwpos120_68 in120_68 sp120_68 202000.000000
Rwpos120_69 in120_69 sp120_69 78000.000000
Rwpos120_70 in120_70 sp120_70 78000.000000
Rwpos120_71 in120_71 sp120_71 202000.000000
Rwpos120_72 in120_72 sp120_72 78000.000000
Rwpos120_73 in120_73 sp120_73 78000.000000
Rwpos120_74 in120_74 sp120_74 78000.000000
Rwpos120_75 in120_75 sp120_75 202000.000000
Rwpos120_76 in120_76 sp120_76 202000.000000
Rwpos120_77 in120_77 sp120_77 202000.000000
Rwpos120_78 in120_78 sp120_78 78000.000000
Rwpos120_79 in120_79 sp120_79 202000.000000
Rwpos120_80 in120_80 sp120_80 78000.000000
Rwpos120_81 in120_81 sp120_81 202000.000000
Rwpos120_82 in120_82 sp120_82 202000.000000
Rwpos120_83 in120_83 sp120_83 78000.000000
Rwpos120_84 in120_84 sp120_84 202000.000000


**********Negative Weighted Array**********

Rwneg1_1 in1_1 sn1_1 202000.000000
Rwneg1_2 in1_2 sn1_2 78000.000000
Rwneg1_3 in1_3 sn1_3 202000.000000
Rwneg1_4 in1_4 sn1_4 78000.000000
Rwneg1_5 in1_5 sn1_5 78000.000000
Rwneg1_6 in1_6 sn1_6 202000.000000
Rwneg1_7 in1_7 sn1_7 202000.000000
Rwneg1_8 in1_8 sn1_8 78000.000000
Rwneg1_9 in1_9 sn1_9 78000.000000
Rwneg1_10 in1_10 sn1_10 202000.000000
Rwneg1_11 in1_11 sn1_11 202000.000000
Rwneg1_12 in1_12 sn1_12 202000.000000
Rwneg1_13 in1_13 sn1_13 78000.000000
Rwneg1_14 in1_14 sn1_14 78000.000000
Rwneg1_15 in1_15 sn1_15 78000.000000
Rwneg1_16 in1_16 sn1_16 78000.000000
Rwneg1_17 in1_17 sn1_17 202000.000000
Rwneg1_18 in1_18 sn1_18 202000.000000
Rwneg1_19 in1_19 sn1_19 78000.000000
Rwneg1_20 in1_20 sn1_20 78000.000000
Rwneg1_21 in1_21 sn1_21 202000.000000
Rwneg1_22 in1_22 sn1_22 78000.000000
Rwneg1_23 in1_23 sn1_23 202000.000000
Rwneg1_24 in1_24 sn1_24 202000.000000
Rwneg1_25 in1_25 sn1_25 202000.000000
Rwneg1_26 in1_26 sn1_26 202000.000000
Rwneg1_27 in1_27 sn1_27 78000.000000
Rwneg1_28 in1_28 sn1_28 78000.000000
Rwneg1_29 in1_29 sn1_29 78000.000000
Rwneg1_30 in1_30 sn1_30 78000.000000
Rwneg1_31 in1_31 sn1_31 202000.000000
Rwneg1_32 in1_32 sn1_32 202000.000000
Rwneg1_33 in1_33 sn1_33 78000.000000
Rwneg1_34 in1_34 sn1_34 78000.000000
Rwneg1_35 in1_35 sn1_35 202000.000000
Rwneg1_36 in1_36 sn1_36 78000.000000
Rwneg1_37 in1_37 sn1_37 78000.000000
Rwneg1_38 in1_38 sn1_38 78000.000000
Rwneg1_39 in1_39 sn1_39 78000.000000
Rwneg1_40 in1_40 sn1_40 78000.000000
Rwneg1_41 in1_41 sn1_41 78000.000000
Rwneg1_42 in1_42 sn1_42 202000.000000
Rwneg1_43 in1_43 sn1_43 202000.000000
Rwneg1_44 in1_44 sn1_44 78000.000000
Rwneg1_45 in1_45 sn1_45 78000.000000
Rwneg1_46 in1_46 sn1_46 78000.000000
Rwneg1_47 in1_47 sn1_47 202000.000000
Rwneg1_48 in1_48 sn1_48 78000.000000
Rwneg1_49 in1_49 sn1_49 78000.000000
Rwneg1_50 in1_50 sn1_50 78000.000000
Rwneg1_51 in1_51 sn1_51 202000.000000
Rwneg1_52 in1_52 sn1_52 78000.000000
Rwneg1_53 in1_53 sn1_53 78000.000000
Rwneg1_54 in1_54 sn1_54 202000.000000
Rwneg1_55 in1_55 sn1_55 202000.000000
Rwneg1_56 in1_56 sn1_56 202000.000000
Rwneg1_57 in1_57 sn1_57 202000.000000
Rwneg1_58 in1_58 sn1_58 78000.000000
Rwneg1_59 in1_59 sn1_59 202000.000000
Rwneg1_60 in1_60 sn1_60 202000.000000
Rwneg1_61 in1_61 sn1_61 78000.000000
Rwneg1_62 in1_62 sn1_62 202000.000000
Rwneg1_63 in1_63 sn1_63 202000.000000
Rwneg1_64 in1_64 sn1_64 202000.000000
Rwneg1_65 in1_65 sn1_65 202000.000000
Rwneg1_66 in1_66 sn1_66 202000.000000
Rwneg1_67 in1_67 sn1_67 78000.000000
Rwneg1_68 in1_68 sn1_68 202000.000000
Rwneg1_69 in1_69 sn1_69 202000.000000
Rwneg1_70 in1_70 sn1_70 78000.000000
Rwneg1_71 in1_71 sn1_71 202000.000000
Rwneg1_72 in1_72 sn1_72 78000.000000
Rwneg1_73 in1_73 sn1_73 202000.000000
Rwneg1_74 in1_74 sn1_74 78000.000000
Rwneg1_75 in1_75 sn1_75 202000.000000
Rwneg1_76 in1_76 sn1_76 78000.000000
Rwneg1_77 in1_77 sn1_77 202000.000000
Rwneg1_78 in1_78 sn1_78 202000.000000
Rwneg1_79 in1_79 sn1_79 202000.000000
Rwneg1_80 in1_80 sn1_80 202000.000000
Rwneg1_81 in1_81 sn1_81 202000.000000
Rwneg1_82 in1_82 sn1_82 78000.000000
Rwneg1_83 in1_83 sn1_83 202000.000000
Rwneg1_84 in1_84 sn1_84 202000.000000
Rwneg2_1 in2_1 sn2_1 202000.000000
Rwneg2_2 in2_2 sn2_2 202000.000000
Rwneg2_3 in2_3 sn2_3 78000.000000
Rwneg2_4 in2_4 sn2_4 202000.000000
Rwneg2_5 in2_5 sn2_5 202000.000000
Rwneg2_6 in2_6 sn2_6 202000.000000
Rwneg2_7 in2_7 sn2_7 78000.000000
Rwneg2_8 in2_8 sn2_8 202000.000000
Rwneg2_9 in2_9 sn2_9 78000.000000
Rwneg2_10 in2_10 sn2_10 202000.000000
Rwneg2_11 in2_11 sn2_11 202000.000000
Rwneg2_12 in2_12 sn2_12 78000.000000
Rwneg2_13 in2_13 sn2_13 202000.000000
Rwneg2_14 in2_14 sn2_14 202000.000000
Rwneg2_15 in2_15 sn2_15 78000.000000
Rwneg2_16 in2_16 sn2_16 78000.000000
Rwneg2_17 in2_17 sn2_17 202000.000000
Rwneg2_18 in2_18 sn2_18 202000.000000
Rwneg2_19 in2_19 sn2_19 78000.000000
Rwneg2_20 in2_20 sn2_20 78000.000000
Rwneg2_21 in2_21 sn2_21 202000.000000
Rwneg2_22 in2_22 sn2_22 202000.000000
Rwneg2_23 in2_23 sn2_23 202000.000000
Rwneg2_24 in2_24 sn2_24 202000.000000
Rwneg2_25 in2_25 sn2_25 78000.000000
Rwneg2_26 in2_26 sn2_26 202000.000000
Rwneg2_27 in2_27 sn2_27 78000.000000
Rwneg2_28 in2_28 sn2_28 78000.000000
Rwneg2_29 in2_29 sn2_29 202000.000000
Rwneg2_30 in2_30 sn2_30 202000.000000
Rwneg2_31 in2_31 sn2_31 78000.000000
Rwneg2_32 in2_32 sn2_32 78000.000000
Rwneg2_33 in2_33 sn2_33 78000.000000
Rwneg2_34 in2_34 sn2_34 78000.000000
Rwneg2_35 in2_35 sn2_35 78000.000000
Rwneg2_36 in2_36 sn2_36 78000.000000
Rwneg2_37 in2_37 sn2_37 78000.000000
Rwneg2_38 in2_38 sn2_38 78000.000000
Rwneg2_39 in2_39 sn2_39 202000.000000
Rwneg2_40 in2_40 sn2_40 78000.000000
Rwneg2_41 in2_41 sn2_41 78000.000000
Rwneg2_42 in2_42 sn2_42 78000.000000
Rwneg2_43 in2_43 sn2_43 202000.000000
Rwneg2_44 in2_44 sn2_44 202000.000000
Rwneg2_45 in2_45 sn2_45 202000.000000
Rwneg2_46 in2_46 sn2_46 78000.000000
Rwneg2_47 in2_47 sn2_47 202000.000000
Rwneg2_48 in2_48 sn2_48 78000.000000
Rwneg2_49 in2_49 sn2_49 78000.000000
Rwneg2_50 in2_50 sn2_50 78000.000000
Rwneg2_51 in2_51 sn2_51 78000.000000
Rwneg2_52 in2_52 sn2_52 78000.000000
Rwneg2_53 in2_53 sn2_53 202000.000000
Rwneg2_54 in2_54 sn2_54 78000.000000
Rwneg2_55 in2_55 sn2_55 202000.000000
Rwneg2_56 in2_56 sn2_56 202000.000000
Rwneg2_57 in2_57 sn2_57 202000.000000
Rwneg2_58 in2_58 sn2_58 202000.000000
Rwneg2_59 in2_59 sn2_59 78000.000000
Rwneg2_60 in2_60 sn2_60 202000.000000
Rwneg2_61 in2_61 sn2_61 202000.000000
Rwneg2_62 in2_62 sn2_62 202000.000000
Rwneg2_63 in2_63 sn2_63 202000.000000
Rwneg2_64 in2_64 sn2_64 78000.000000
Rwneg2_65 in2_65 sn2_65 202000.000000
Rwneg2_66 in2_66 sn2_66 78000.000000
Rwneg2_67 in2_67 sn2_67 78000.000000
Rwneg2_68 in2_68 sn2_68 202000.000000
Rwneg2_69 in2_69 sn2_69 202000.000000
Rwneg2_70 in2_70 sn2_70 202000.000000
Rwneg2_71 in2_71 sn2_71 202000.000000
Rwneg2_72 in2_72 sn2_72 202000.000000
Rwneg2_73 in2_73 sn2_73 202000.000000
Rwneg2_74 in2_74 sn2_74 202000.000000
Rwneg2_75 in2_75 sn2_75 78000.000000
Rwneg2_76 in2_76 sn2_76 78000.000000
Rwneg2_77 in2_77 sn2_77 78000.000000
Rwneg2_78 in2_78 sn2_78 78000.000000
Rwneg2_79 in2_79 sn2_79 202000.000000
Rwneg2_80 in2_80 sn2_80 202000.000000
Rwneg2_81 in2_81 sn2_81 202000.000000
Rwneg2_82 in2_82 sn2_82 202000.000000
Rwneg2_83 in2_83 sn2_83 202000.000000
Rwneg2_84 in2_84 sn2_84 202000.000000
Rwneg3_1 in3_1 sn3_1 78000.000000
Rwneg3_2 in3_2 sn3_2 78000.000000
Rwneg3_3 in3_3 sn3_3 78000.000000
Rwneg3_4 in3_4 sn3_4 202000.000000
Rwneg3_5 in3_5 sn3_5 78000.000000
Rwneg3_6 in3_6 sn3_6 202000.000000
Rwneg3_7 in3_7 sn3_7 202000.000000
Rwneg3_8 in3_8 sn3_8 78000.000000
Rwneg3_9 in3_9 sn3_9 78000.000000
Rwneg3_10 in3_10 sn3_10 202000.000000
Rwneg3_11 in3_11 sn3_11 202000.000000
Rwneg3_12 in3_12 sn3_12 202000.000000
Rwneg3_13 in3_13 sn3_13 202000.000000
Rwneg3_14 in3_14 sn3_14 202000.000000
Rwneg3_15 in3_15 sn3_15 202000.000000
Rwneg3_16 in3_16 sn3_16 202000.000000
Rwneg3_17 in3_17 sn3_17 78000.000000
Rwneg3_18 in3_18 sn3_18 202000.000000
Rwneg3_19 in3_19 sn3_19 202000.000000
Rwneg3_20 in3_20 sn3_20 202000.000000
Rwneg3_21 in3_21 sn3_21 78000.000000
Rwneg3_22 in3_22 sn3_22 78000.000000
Rwneg3_23 in3_23 sn3_23 78000.000000
Rwneg3_24 in3_24 sn3_24 202000.000000
Rwneg3_25 in3_25 sn3_25 78000.000000
Rwneg3_26 in3_26 sn3_26 202000.000000
Rwneg3_27 in3_27 sn3_27 202000.000000
Rwneg3_28 in3_28 sn3_28 202000.000000
Rwneg3_29 in3_29 sn3_29 78000.000000
Rwneg3_30 in3_30 sn3_30 78000.000000
Rwneg3_31 in3_31 sn3_31 78000.000000
Rwneg3_32 in3_32 sn3_32 202000.000000
Rwneg3_33 in3_33 sn3_33 78000.000000
Rwneg3_34 in3_34 sn3_34 202000.000000
Rwneg3_35 in3_35 sn3_35 78000.000000
Rwneg3_36 in3_36 sn3_36 202000.000000
Rwneg3_37 in3_37 sn3_37 202000.000000
Rwneg3_38 in3_38 sn3_38 202000.000000
Rwneg3_39 in3_39 sn3_39 202000.000000
Rwneg3_40 in3_40 sn3_40 202000.000000
Rwneg3_41 in3_41 sn3_41 78000.000000
Rwneg3_42 in3_42 sn3_42 78000.000000
Rwneg3_43 in3_43 sn3_43 202000.000000
Rwneg3_44 in3_44 sn3_44 78000.000000
Rwneg3_45 in3_45 sn3_45 202000.000000
Rwneg3_46 in3_46 sn3_46 202000.000000
Rwneg3_47 in3_47 sn3_47 202000.000000
Rwneg3_48 in3_48 sn3_48 78000.000000
Rwneg3_49 in3_49 sn3_49 202000.000000
Rwneg3_50 in3_50 sn3_50 202000.000000
Rwneg3_51 in3_51 sn3_51 202000.000000
Rwneg3_52 in3_52 sn3_52 202000.000000
Rwneg3_53 in3_53 sn3_53 78000.000000
Rwneg3_54 in3_54 sn3_54 202000.000000
Rwneg3_55 in3_55 sn3_55 78000.000000
Rwneg3_56 in3_56 sn3_56 202000.000000
Rwneg3_57 in3_57 sn3_57 202000.000000
Rwneg3_58 in3_58 sn3_58 78000.000000
Rwneg3_59 in3_59 sn3_59 202000.000000
Rwneg3_60 in3_60 sn3_60 202000.000000
Rwneg3_61 in3_61 sn3_61 78000.000000
Rwneg3_62 in3_62 sn3_62 78000.000000
Rwneg3_63 in3_63 sn3_63 202000.000000
Rwneg3_64 in3_64 sn3_64 78000.000000
Rwneg3_65 in3_65 sn3_65 78000.000000
Rwneg3_66 in3_66 sn3_66 78000.000000
Rwneg3_67 in3_67 sn3_67 202000.000000
Rwneg3_68 in3_68 sn3_68 202000.000000
Rwneg3_69 in3_69 sn3_69 202000.000000
Rwneg3_70 in3_70 sn3_70 78000.000000
Rwneg3_71 in3_71 sn3_71 78000.000000
Rwneg3_72 in3_72 sn3_72 202000.000000
Rwneg3_73 in3_73 sn3_73 78000.000000
Rwneg3_74 in3_74 sn3_74 78000.000000
Rwneg3_75 in3_75 sn3_75 202000.000000
Rwneg3_76 in3_76 sn3_76 202000.000000
Rwneg3_77 in3_77 sn3_77 202000.000000
Rwneg3_78 in3_78 sn3_78 202000.000000
Rwneg3_79 in3_79 sn3_79 202000.000000
Rwneg3_80 in3_80 sn3_80 78000.000000
Rwneg3_81 in3_81 sn3_81 78000.000000
Rwneg3_82 in3_82 sn3_82 202000.000000
Rwneg3_83 in3_83 sn3_83 78000.000000
Rwneg3_84 in3_84 sn3_84 78000.000000
Rwneg4_1 in4_1 sn4_1 78000.000000
Rwneg4_2 in4_2 sn4_2 78000.000000
Rwneg4_3 in4_3 sn4_3 78000.000000
Rwneg4_4 in4_4 sn4_4 202000.000000
Rwneg4_5 in4_5 sn4_5 202000.000000
Rwneg4_6 in4_6 sn4_6 202000.000000
Rwneg4_7 in4_7 sn4_7 202000.000000
Rwneg4_8 in4_8 sn4_8 78000.000000
Rwneg4_9 in4_9 sn4_9 202000.000000
Rwneg4_10 in4_10 sn4_10 78000.000000
Rwneg4_11 in4_11 sn4_11 202000.000000
Rwneg4_12 in4_12 sn4_12 78000.000000
Rwneg4_13 in4_13 sn4_13 202000.000000
Rwneg4_14 in4_14 sn4_14 202000.000000
Rwneg4_15 in4_15 sn4_15 202000.000000
Rwneg4_16 in4_16 sn4_16 78000.000000
Rwneg4_17 in4_17 sn4_17 202000.000000
Rwneg4_18 in4_18 sn4_18 202000.000000
Rwneg4_19 in4_19 sn4_19 78000.000000
Rwneg4_20 in4_20 sn4_20 78000.000000
Rwneg4_21 in4_21 sn4_21 202000.000000
Rwneg4_22 in4_22 sn4_22 78000.000000
Rwneg4_23 in4_23 sn4_23 202000.000000
Rwneg4_24 in4_24 sn4_24 202000.000000
Rwneg4_25 in4_25 sn4_25 202000.000000
Rwneg4_26 in4_26 sn4_26 202000.000000
Rwneg4_27 in4_27 sn4_27 202000.000000
Rwneg4_28 in4_28 sn4_28 202000.000000
Rwneg4_29 in4_29 sn4_29 78000.000000
Rwneg4_30 in4_30 sn4_30 202000.000000
Rwneg4_31 in4_31 sn4_31 202000.000000
Rwneg4_32 in4_32 sn4_32 202000.000000
Rwneg4_33 in4_33 sn4_33 78000.000000
Rwneg4_34 in4_34 sn4_34 202000.000000
Rwneg4_35 in4_35 sn4_35 202000.000000
Rwneg4_36 in4_36 sn4_36 78000.000000
Rwneg4_37 in4_37 sn4_37 202000.000000
Rwneg4_38 in4_38 sn4_38 78000.000000
Rwneg4_39 in4_39 sn4_39 202000.000000
Rwneg4_40 in4_40 sn4_40 78000.000000
Rwneg4_41 in4_41 sn4_41 78000.000000
Rwneg4_42 in4_42 sn4_42 202000.000000
Rwneg4_43 in4_43 sn4_43 202000.000000
Rwneg4_44 in4_44 sn4_44 78000.000000
Rwneg4_45 in4_45 sn4_45 78000.000000
Rwneg4_46 in4_46 sn4_46 202000.000000
Rwneg4_47 in4_47 sn4_47 202000.000000
Rwneg4_48 in4_48 sn4_48 78000.000000
Rwneg4_49 in4_49 sn4_49 78000.000000
Rwneg4_50 in4_50 sn4_50 202000.000000
Rwneg4_51 in4_51 sn4_51 202000.000000
Rwneg4_52 in4_52 sn4_52 202000.000000
Rwneg4_53 in4_53 sn4_53 78000.000000
Rwneg4_54 in4_54 sn4_54 202000.000000
Rwneg4_55 in4_55 sn4_55 78000.000000
Rwneg4_56 in4_56 sn4_56 78000.000000
Rwneg4_57 in4_57 sn4_57 78000.000000
Rwneg4_58 in4_58 sn4_58 78000.000000
Rwneg4_59 in4_59 sn4_59 78000.000000
Rwneg4_60 in4_60 sn4_60 202000.000000
Rwneg4_61 in4_61 sn4_61 78000.000000
Rwneg4_62 in4_62 sn4_62 202000.000000
Rwneg4_63 in4_63 sn4_63 78000.000000
Rwneg4_64 in4_64 sn4_64 78000.000000
Rwneg4_65 in4_65 sn4_65 78000.000000
Rwneg4_66 in4_66 sn4_66 78000.000000
Rwneg4_67 in4_67 sn4_67 78000.000000
Rwneg4_68 in4_68 sn4_68 78000.000000
Rwneg4_69 in4_69 sn4_69 78000.000000
Rwneg4_70 in4_70 sn4_70 78000.000000
Rwneg4_71 in4_71 sn4_71 78000.000000
Rwneg4_72 in4_72 sn4_72 78000.000000
Rwneg4_73 in4_73 sn4_73 78000.000000
Rwneg4_74 in4_74 sn4_74 78000.000000
Rwneg4_75 in4_75 sn4_75 78000.000000
Rwneg4_76 in4_76 sn4_76 78000.000000
Rwneg4_77 in4_77 sn4_77 202000.000000
Rwneg4_78 in4_78 sn4_78 202000.000000
Rwneg4_79 in4_79 sn4_79 78000.000000
Rwneg4_80 in4_80 sn4_80 202000.000000
Rwneg4_81 in4_81 sn4_81 202000.000000
Rwneg4_82 in4_82 sn4_82 78000.000000
Rwneg4_83 in4_83 sn4_83 78000.000000
Rwneg4_84 in4_84 sn4_84 78000.000000
Rwneg5_1 in5_1 sn5_1 202000.000000
Rwneg5_2 in5_2 sn5_2 202000.000000
Rwneg5_3 in5_3 sn5_3 78000.000000
Rwneg5_4 in5_4 sn5_4 202000.000000
Rwneg5_5 in5_5 sn5_5 202000.000000
Rwneg5_6 in5_6 sn5_6 202000.000000
Rwneg5_7 in5_7 sn5_7 78000.000000
Rwneg5_8 in5_8 sn5_8 202000.000000
Rwneg5_9 in5_9 sn5_9 202000.000000
Rwneg5_10 in5_10 sn5_10 202000.000000
Rwneg5_11 in5_11 sn5_11 202000.000000
Rwneg5_12 in5_12 sn5_12 202000.000000
Rwneg5_13 in5_13 sn5_13 202000.000000
Rwneg5_14 in5_14 sn5_14 78000.000000
Rwneg5_15 in5_15 sn5_15 202000.000000
Rwneg5_16 in5_16 sn5_16 202000.000000
Rwneg5_17 in5_17 sn5_17 78000.000000
Rwneg5_18 in5_18 sn5_18 202000.000000
Rwneg5_19 in5_19 sn5_19 202000.000000
Rwneg5_20 in5_20 sn5_20 78000.000000
Rwneg5_21 in5_21 sn5_21 78000.000000
Rwneg5_22 in5_22 sn5_22 78000.000000
Rwneg5_23 in5_23 sn5_23 78000.000000
Rwneg5_24 in5_24 sn5_24 202000.000000
Rwneg5_25 in5_25 sn5_25 78000.000000
Rwneg5_26 in5_26 sn5_26 202000.000000
Rwneg5_27 in5_27 sn5_27 202000.000000
Rwneg5_28 in5_28 sn5_28 202000.000000
Rwneg5_29 in5_29 sn5_29 202000.000000
Rwneg5_30 in5_30 sn5_30 202000.000000
Rwneg5_31 in5_31 sn5_31 202000.000000
Rwneg5_32 in5_32 sn5_32 78000.000000
Rwneg5_33 in5_33 sn5_33 78000.000000
Rwneg5_34 in5_34 sn5_34 78000.000000
Rwneg5_35 in5_35 sn5_35 78000.000000
Rwneg5_36 in5_36 sn5_36 78000.000000
Rwneg5_37 in5_37 sn5_37 78000.000000
Rwneg5_38 in5_38 sn5_38 202000.000000
Rwneg5_39 in5_39 sn5_39 78000.000000
Rwneg5_40 in5_40 sn5_40 202000.000000
Rwneg5_41 in5_41 sn5_41 202000.000000
Rwneg5_42 in5_42 sn5_42 202000.000000
Rwneg5_43 in5_43 sn5_43 202000.000000
Rwneg5_44 in5_44 sn5_44 202000.000000
Rwneg5_45 in5_45 sn5_45 78000.000000
Rwneg5_46 in5_46 sn5_46 78000.000000
Rwneg5_47 in5_47 sn5_47 78000.000000
Rwneg5_48 in5_48 sn5_48 78000.000000
Rwneg5_49 in5_49 sn5_49 202000.000000
Rwneg5_50 in5_50 sn5_50 78000.000000
Rwneg5_51 in5_51 sn5_51 202000.000000
Rwneg5_52 in5_52 sn5_52 202000.000000
Rwneg5_53 in5_53 sn5_53 78000.000000
Rwneg5_54 in5_54 sn5_54 202000.000000
Rwneg5_55 in5_55 sn5_55 202000.000000
Rwneg5_56 in5_56 sn5_56 78000.000000
Rwneg5_57 in5_57 sn5_57 78000.000000
Rwneg5_58 in5_58 sn5_58 202000.000000
Rwneg5_59 in5_59 sn5_59 78000.000000
Rwneg5_60 in5_60 sn5_60 202000.000000
Rwneg5_61 in5_61 sn5_61 78000.000000
Rwneg5_62 in5_62 sn5_62 202000.000000
Rwneg5_63 in5_63 sn5_63 78000.000000
Rwneg5_64 in5_64 sn5_64 78000.000000
Rwneg5_65 in5_65 sn5_65 78000.000000
Rwneg5_66 in5_66 sn5_66 202000.000000
Rwneg5_67 in5_67 sn5_67 78000.000000
Rwneg5_68 in5_68 sn5_68 202000.000000
Rwneg5_69 in5_69 sn5_69 78000.000000
Rwneg5_70 in5_70 sn5_70 202000.000000
Rwneg5_71 in5_71 sn5_71 78000.000000
Rwneg5_72 in5_72 sn5_72 78000.000000
Rwneg5_73 in5_73 sn5_73 202000.000000
Rwneg5_74 in5_74 sn5_74 78000.000000
Rwneg5_75 in5_75 sn5_75 78000.000000
Rwneg5_76 in5_76 sn5_76 202000.000000
Rwneg5_77 in5_77 sn5_77 78000.000000
Rwneg5_78 in5_78 sn5_78 202000.000000
Rwneg5_79 in5_79 sn5_79 78000.000000
Rwneg5_80 in5_80 sn5_80 78000.000000
Rwneg5_81 in5_81 sn5_81 78000.000000
Rwneg5_82 in5_82 sn5_82 202000.000000
Rwneg5_83 in5_83 sn5_83 78000.000000
Rwneg5_84 in5_84 sn5_84 202000.000000
Rwneg6_1 in6_1 sn6_1 78000.000000
Rwneg6_2 in6_2 sn6_2 202000.000000
Rwneg6_3 in6_3 sn6_3 78000.000000
Rwneg6_4 in6_4 sn6_4 202000.000000
Rwneg6_5 in6_5 sn6_5 78000.000000
Rwneg6_6 in6_6 sn6_6 202000.000000
Rwneg6_7 in6_7 sn6_7 78000.000000
Rwneg6_8 in6_8 sn6_8 78000.000000
Rwneg6_9 in6_9 sn6_9 202000.000000
Rwneg6_10 in6_10 sn6_10 202000.000000
Rwneg6_11 in6_11 sn6_11 78000.000000
Rwneg6_12 in6_12 sn6_12 202000.000000
Rwneg6_13 in6_13 sn6_13 78000.000000
Rwneg6_14 in6_14 sn6_14 78000.000000
Rwneg6_15 in6_15 sn6_15 78000.000000
Rwneg6_16 in6_16 sn6_16 202000.000000
Rwneg6_17 in6_17 sn6_17 78000.000000
Rwneg6_18 in6_18 sn6_18 78000.000000
Rwneg6_19 in6_19 sn6_19 202000.000000
Rwneg6_20 in6_20 sn6_20 202000.000000
Rwneg6_21 in6_21 sn6_21 78000.000000
Rwneg6_22 in6_22 sn6_22 78000.000000
Rwneg6_23 in6_23 sn6_23 78000.000000
Rwneg6_24 in6_24 sn6_24 78000.000000
Rwneg6_25 in6_25 sn6_25 78000.000000
Rwneg6_26 in6_26 sn6_26 78000.000000
Rwneg6_27 in6_27 sn6_27 78000.000000
Rwneg6_28 in6_28 sn6_28 202000.000000
Rwneg6_29 in6_29 sn6_29 202000.000000
Rwneg6_30 in6_30 sn6_30 202000.000000
Rwneg6_31 in6_31 sn6_31 78000.000000
Rwneg6_32 in6_32 sn6_32 78000.000000
Rwneg6_33 in6_33 sn6_33 202000.000000
Rwneg6_34 in6_34 sn6_34 202000.000000
Rwneg6_35 in6_35 sn6_35 202000.000000
Rwneg6_36 in6_36 sn6_36 78000.000000
Rwneg6_37 in6_37 sn6_37 78000.000000
Rwneg6_38 in6_38 sn6_38 202000.000000
Rwneg6_39 in6_39 sn6_39 78000.000000
Rwneg6_40 in6_40 sn6_40 202000.000000
Rwneg6_41 in6_41 sn6_41 78000.000000
Rwneg6_42 in6_42 sn6_42 78000.000000
Rwneg6_43 in6_43 sn6_43 202000.000000
Rwneg6_44 in6_44 sn6_44 78000.000000
Rwneg6_45 in6_45 sn6_45 202000.000000
Rwneg6_46 in6_46 sn6_46 78000.000000
Rwneg6_47 in6_47 sn6_47 202000.000000
Rwneg6_48 in6_48 sn6_48 78000.000000
Rwneg6_49 in6_49 sn6_49 202000.000000
Rwneg6_50 in6_50 sn6_50 78000.000000
Rwneg6_51 in6_51 sn6_51 78000.000000
Rwneg6_52 in6_52 sn6_52 202000.000000
Rwneg6_53 in6_53 sn6_53 202000.000000
Rwneg6_54 in6_54 sn6_54 78000.000000
Rwneg6_55 in6_55 sn6_55 202000.000000
Rwneg6_56 in6_56 sn6_56 78000.000000
Rwneg6_57 in6_57 sn6_57 78000.000000
Rwneg6_58 in6_58 sn6_58 78000.000000
Rwneg6_59 in6_59 sn6_59 78000.000000
Rwneg6_60 in6_60 sn6_60 202000.000000
Rwneg6_61 in6_61 sn6_61 202000.000000
Rwneg6_62 in6_62 sn6_62 78000.000000
Rwneg6_63 in6_63 sn6_63 202000.000000
Rwneg6_64 in6_64 sn6_64 78000.000000
Rwneg6_65 in6_65 sn6_65 202000.000000
Rwneg6_66 in6_66 sn6_66 78000.000000
Rwneg6_67 in6_67 sn6_67 202000.000000
Rwneg6_68 in6_68 sn6_68 78000.000000
Rwneg6_69 in6_69 sn6_69 78000.000000
Rwneg6_70 in6_70 sn6_70 202000.000000
Rwneg6_71 in6_71 sn6_71 78000.000000
Rwneg6_72 in6_72 sn6_72 202000.000000
Rwneg6_73 in6_73 sn6_73 78000.000000
Rwneg6_74 in6_74 sn6_74 78000.000000
Rwneg6_75 in6_75 sn6_75 202000.000000
Rwneg6_76 in6_76 sn6_76 202000.000000
Rwneg6_77 in6_77 sn6_77 202000.000000
Rwneg6_78 in6_78 sn6_78 202000.000000
Rwneg6_79 in6_79 sn6_79 78000.000000
Rwneg6_80 in6_80 sn6_80 78000.000000
Rwneg6_81 in6_81 sn6_81 78000.000000
Rwneg6_82 in6_82 sn6_82 78000.000000
Rwneg6_83 in6_83 sn6_83 78000.000000
Rwneg6_84 in6_84 sn6_84 78000.000000
Rwneg7_1 in7_1 sn7_1 202000.000000
Rwneg7_2 in7_2 sn7_2 78000.000000
Rwneg7_3 in7_3 sn7_3 78000.000000
Rwneg7_4 in7_4 sn7_4 78000.000000
Rwneg7_5 in7_5 sn7_5 202000.000000
Rwneg7_6 in7_6 sn7_6 202000.000000
Rwneg7_7 in7_7 sn7_7 202000.000000
Rwneg7_8 in7_8 sn7_8 78000.000000
Rwneg7_9 in7_9 sn7_9 202000.000000
Rwneg7_10 in7_10 sn7_10 202000.000000
Rwneg7_11 in7_11 sn7_11 78000.000000
Rwneg7_12 in7_12 sn7_12 202000.000000
Rwneg7_13 in7_13 sn7_13 78000.000000
Rwneg7_14 in7_14 sn7_14 202000.000000
Rwneg7_15 in7_15 sn7_15 78000.000000
Rwneg7_16 in7_16 sn7_16 78000.000000
Rwneg7_17 in7_17 sn7_17 202000.000000
Rwneg7_18 in7_18 sn7_18 202000.000000
Rwneg7_19 in7_19 sn7_19 78000.000000
Rwneg7_20 in7_20 sn7_20 78000.000000
Rwneg7_21 in7_21 sn7_21 78000.000000
Rwneg7_22 in7_22 sn7_22 78000.000000
Rwneg7_23 in7_23 sn7_23 78000.000000
Rwneg7_24 in7_24 sn7_24 202000.000000
Rwneg7_25 in7_25 sn7_25 202000.000000
Rwneg7_26 in7_26 sn7_26 78000.000000
Rwneg7_27 in7_27 sn7_27 202000.000000
Rwneg7_28 in7_28 sn7_28 202000.000000
Rwneg7_29 in7_29 sn7_29 202000.000000
Rwneg7_30 in7_30 sn7_30 202000.000000
Rwneg7_31 in7_31 sn7_31 78000.000000
Rwneg7_32 in7_32 sn7_32 202000.000000
Rwneg7_33 in7_33 sn7_33 78000.000000
Rwneg7_34 in7_34 sn7_34 202000.000000
Rwneg7_35 in7_35 sn7_35 78000.000000
Rwneg7_36 in7_36 sn7_36 202000.000000
Rwneg7_37 in7_37 sn7_37 78000.000000
Rwneg7_38 in7_38 sn7_38 202000.000000
Rwneg7_39 in7_39 sn7_39 202000.000000
Rwneg7_40 in7_40 sn7_40 78000.000000
Rwneg7_41 in7_41 sn7_41 78000.000000
Rwneg7_42 in7_42 sn7_42 202000.000000
Rwneg7_43 in7_43 sn7_43 202000.000000
Rwneg7_44 in7_44 sn7_44 202000.000000
Rwneg7_45 in7_45 sn7_45 78000.000000
Rwneg7_46 in7_46 sn7_46 202000.000000
Rwneg7_47 in7_47 sn7_47 202000.000000
Rwneg7_48 in7_48 sn7_48 78000.000000
Rwneg7_49 in7_49 sn7_49 202000.000000
Rwneg7_50 in7_50 sn7_50 78000.000000
Rwneg7_51 in7_51 sn7_51 78000.000000
Rwneg7_52 in7_52 sn7_52 202000.000000
Rwneg7_53 in7_53 sn7_53 202000.000000
Rwneg7_54 in7_54 sn7_54 78000.000000
Rwneg7_55 in7_55 sn7_55 78000.000000
Rwneg7_56 in7_56 sn7_56 78000.000000
Rwneg7_57 in7_57 sn7_57 78000.000000
Rwneg7_58 in7_58 sn7_58 78000.000000
Rwneg7_59 in7_59 sn7_59 78000.000000
Rwneg7_60 in7_60 sn7_60 202000.000000
Rwneg7_61 in7_61 sn7_61 78000.000000
Rwneg7_62 in7_62 sn7_62 202000.000000
Rwneg7_63 in7_63 sn7_63 202000.000000
Rwneg7_64 in7_64 sn7_64 202000.000000
Rwneg7_65 in7_65 sn7_65 202000.000000
Rwneg7_66 in7_66 sn7_66 202000.000000
Rwneg7_67 in7_67 sn7_67 202000.000000
Rwneg7_68 in7_68 sn7_68 202000.000000
Rwneg7_69 in7_69 sn7_69 202000.000000
Rwneg7_70 in7_70 sn7_70 202000.000000
Rwneg7_71 in7_71 sn7_71 202000.000000
Rwneg7_72 in7_72 sn7_72 202000.000000
Rwneg7_73 in7_73 sn7_73 78000.000000
Rwneg7_74 in7_74 sn7_74 202000.000000
Rwneg7_75 in7_75 sn7_75 78000.000000
Rwneg7_76 in7_76 sn7_76 202000.000000
Rwneg7_77 in7_77 sn7_77 202000.000000
Rwneg7_78 in7_78 sn7_78 202000.000000
Rwneg7_79 in7_79 sn7_79 202000.000000
Rwneg7_80 in7_80 sn7_80 78000.000000
Rwneg7_81 in7_81 sn7_81 78000.000000
Rwneg7_82 in7_82 sn7_82 202000.000000
Rwneg7_83 in7_83 sn7_83 78000.000000
Rwneg7_84 in7_84 sn7_84 78000.000000
Rwneg8_1 in8_1 sn8_1 78000.000000
Rwneg8_2 in8_2 sn8_2 202000.000000
Rwneg8_3 in8_3 sn8_3 202000.000000
Rwneg8_4 in8_4 sn8_4 78000.000000
Rwneg8_5 in8_5 sn8_5 78000.000000
Rwneg8_6 in8_6 sn8_6 202000.000000
Rwneg8_7 in8_7 sn8_7 202000.000000
Rwneg8_8 in8_8 sn8_8 78000.000000
Rwneg8_9 in8_9 sn8_9 78000.000000
Rwneg8_10 in8_10 sn8_10 78000.000000
Rwneg8_11 in8_11 sn8_11 78000.000000
Rwneg8_12 in8_12 sn8_12 78000.000000
Rwneg8_13 in8_13 sn8_13 78000.000000
Rwneg8_14 in8_14 sn8_14 202000.000000
Rwneg8_15 in8_15 sn8_15 78000.000000
Rwneg8_16 in8_16 sn8_16 78000.000000
Rwneg8_17 in8_17 sn8_17 202000.000000
Rwneg8_18 in8_18 sn8_18 78000.000000
Rwneg8_19 in8_19 sn8_19 78000.000000
Rwneg8_20 in8_20 sn8_20 78000.000000
Rwneg8_21 in8_21 sn8_21 78000.000000
Rwneg8_22 in8_22 sn8_22 78000.000000
Rwneg8_23 in8_23 sn8_23 202000.000000
Rwneg8_24 in8_24 sn8_24 202000.000000
Rwneg8_25 in8_25 sn8_25 78000.000000
Rwneg8_26 in8_26 sn8_26 202000.000000
Rwneg8_27 in8_27 sn8_27 78000.000000
Rwneg8_28 in8_28 sn8_28 78000.000000
Rwneg8_29 in8_29 sn8_29 78000.000000
Rwneg8_30 in8_30 sn8_30 202000.000000
Rwneg8_31 in8_31 sn8_31 202000.000000
Rwneg8_32 in8_32 sn8_32 78000.000000
Rwneg8_33 in8_33 sn8_33 202000.000000
Rwneg8_34 in8_34 sn8_34 78000.000000
Rwneg8_35 in8_35 sn8_35 78000.000000
Rwneg8_36 in8_36 sn8_36 78000.000000
Rwneg8_37 in8_37 sn8_37 202000.000000
Rwneg8_38 in8_38 sn8_38 78000.000000
Rwneg8_39 in8_39 sn8_39 78000.000000
Rwneg8_40 in8_40 sn8_40 202000.000000
Rwneg8_41 in8_41 sn8_41 202000.000000
Rwneg8_42 in8_42 sn8_42 202000.000000
Rwneg8_43 in8_43 sn8_43 202000.000000
Rwneg8_44 in8_44 sn8_44 202000.000000
Rwneg8_45 in8_45 sn8_45 78000.000000
Rwneg8_46 in8_46 sn8_46 202000.000000
Rwneg8_47 in8_47 sn8_47 202000.000000
Rwneg8_48 in8_48 sn8_48 78000.000000
Rwneg8_49 in8_49 sn8_49 202000.000000
Rwneg8_50 in8_50 sn8_50 78000.000000
Rwneg8_51 in8_51 sn8_51 202000.000000
Rwneg8_52 in8_52 sn8_52 78000.000000
Rwneg8_53 in8_53 sn8_53 78000.000000
Rwneg8_54 in8_54 sn8_54 78000.000000
Rwneg8_55 in8_55 sn8_55 78000.000000
Rwneg8_56 in8_56 sn8_56 78000.000000
Rwneg8_57 in8_57 sn8_57 202000.000000
Rwneg8_58 in8_58 sn8_58 202000.000000
Rwneg8_59 in8_59 sn8_59 202000.000000
Rwneg8_60 in8_60 sn8_60 202000.000000
Rwneg8_61 in8_61 sn8_61 202000.000000
Rwneg8_62 in8_62 sn8_62 78000.000000
Rwneg8_63 in8_63 sn8_63 78000.000000
Rwneg8_64 in8_64 sn8_64 78000.000000
Rwneg8_65 in8_65 sn8_65 202000.000000
Rwneg8_66 in8_66 sn8_66 78000.000000
Rwneg8_67 in8_67 sn8_67 202000.000000
Rwneg8_68 in8_68 sn8_68 78000.000000
Rwneg8_69 in8_69 sn8_69 202000.000000
Rwneg8_70 in8_70 sn8_70 78000.000000
Rwneg8_71 in8_71 sn8_71 78000.000000
Rwneg8_72 in8_72 sn8_72 202000.000000
Rwneg8_73 in8_73 sn8_73 202000.000000
Rwneg8_74 in8_74 sn8_74 78000.000000
Rwneg8_75 in8_75 sn8_75 202000.000000
Rwneg8_76 in8_76 sn8_76 78000.000000
Rwneg8_77 in8_77 sn8_77 202000.000000
Rwneg8_78 in8_78 sn8_78 78000.000000
Rwneg8_79 in8_79 sn8_79 202000.000000
Rwneg8_80 in8_80 sn8_80 78000.000000
Rwneg8_81 in8_81 sn8_81 202000.000000
Rwneg8_82 in8_82 sn8_82 78000.000000
Rwneg8_83 in8_83 sn8_83 202000.000000
Rwneg8_84 in8_84 sn8_84 78000.000000
Rwneg9_1 in9_1 sn9_1 202000.000000
Rwneg9_2 in9_2 sn9_2 202000.000000
Rwneg9_3 in9_3 sn9_3 202000.000000
Rwneg9_4 in9_4 sn9_4 202000.000000
Rwneg9_5 in9_5 sn9_5 78000.000000
Rwneg9_6 in9_6 sn9_6 202000.000000
Rwneg9_7 in9_7 sn9_7 202000.000000
Rwneg9_8 in9_8 sn9_8 78000.000000
Rwneg9_9 in9_9 sn9_9 202000.000000
Rwneg9_10 in9_10 sn9_10 202000.000000
Rwneg9_11 in9_11 sn9_11 202000.000000
Rwneg9_12 in9_12 sn9_12 202000.000000
Rwneg9_13 in9_13 sn9_13 78000.000000
Rwneg9_14 in9_14 sn9_14 78000.000000
Rwneg9_15 in9_15 sn9_15 202000.000000
Rwneg9_16 in9_16 sn9_16 78000.000000
Rwneg9_17 in9_17 sn9_17 78000.000000
Rwneg9_18 in9_18 sn9_18 78000.000000
Rwneg9_19 in9_19 sn9_19 78000.000000
Rwneg9_20 in9_20 sn9_20 202000.000000
Rwneg9_21 in9_21 sn9_21 202000.000000
Rwneg9_22 in9_22 sn9_22 202000.000000
Rwneg9_23 in9_23 sn9_23 78000.000000
Rwneg9_24 in9_24 sn9_24 202000.000000
Rwneg9_25 in9_25 sn9_25 202000.000000
Rwneg9_26 in9_26 sn9_26 202000.000000
Rwneg9_27 in9_27 sn9_27 78000.000000
Rwneg9_28 in9_28 sn9_28 78000.000000
Rwneg9_29 in9_29 sn9_29 78000.000000
Rwneg9_30 in9_30 sn9_30 202000.000000
Rwneg9_31 in9_31 sn9_31 202000.000000
Rwneg9_32 in9_32 sn9_32 202000.000000
Rwneg9_33 in9_33 sn9_33 202000.000000
Rwneg9_34 in9_34 sn9_34 78000.000000
Rwneg9_35 in9_35 sn9_35 202000.000000
Rwneg9_36 in9_36 sn9_36 202000.000000
Rwneg9_37 in9_37 sn9_37 202000.000000
Rwneg9_38 in9_38 sn9_38 202000.000000
Rwneg9_39 in9_39 sn9_39 78000.000000
Rwneg9_40 in9_40 sn9_40 78000.000000
Rwneg9_41 in9_41 sn9_41 202000.000000
Rwneg9_42 in9_42 sn9_42 202000.000000
Rwneg9_43 in9_43 sn9_43 202000.000000
Rwneg9_44 in9_44 sn9_44 78000.000000
Rwneg9_45 in9_45 sn9_45 202000.000000
Rwneg9_46 in9_46 sn9_46 202000.000000
Rwneg9_47 in9_47 sn9_47 78000.000000
Rwneg9_48 in9_48 sn9_48 202000.000000
Rwneg9_49 in9_49 sn9_49 202000.000000
Rwneg9_50 in9_50 sn9_50 202000.000000
Rwneg9_51 in9_51 sn9_51 78000.000000
Rwneg9_52 in9_52 sn9_52 202000.000000
Rwneg9_53 in9_53 sn9_53 202000.000000
Rwneg9_54 in9_54 sn9_54 78000.000000
Rwneg9_55 in9_55 sn9_55 78000.000000
Rwneg9_56 in9_56 sn9_56 202000.000000
Rwneg9_57 in9_57 sn9_57 202000.000000
Rwneg9_58 in9_58 sn9_58 78000.000000
Rwneg9_59 in9_59 sn9_59 202000.000000
Rwneg9_60 in9_60 sn9_60 202000.000000
Rwneg9_61 in9_61 sn9_61 202000.000000
Rwneg9_62 in9_62 sn9_62 78000.000000
Rwneg9_63 in9_63 sn9_63 202000.000000
Rwneg9_64 in9_64 sn9_64 78000.000000
Rwneg9_65 in9_65 sn9_65 202000.000000
Rwneg9_66 in9_66 sn9_66 202000.000000
Rwneg9_67 in9_67 sn9_67 78000.000000
Rwneg9_68 in9_68 sn9_68 78000.000000
Rwneg9_69 in9_69 sn9_69 78000.000000
Rwneg9_70 in9_70 sn9_70 202000.000000
Rwneg9_71 in9_71 sn9_71 202000.000000
Rwneg9_72 in9_72 sn9_72 202000.000000
Rwneg9_73 in9_73 sn9_73 202000.000000
Rwneg9_74 in9_74 sn9_74 202000.000000
Rwneg9_75 in9_75 sn9_75 202000.000000
Rwneg9_76 in9_76 sn9_76 202000.000000
Rwneg9_77 in9_77 sn9_77 78000.000000
Rwneg9_78 in9_78 sn9_78 202000.000000
Rwneg9_79 in9_79 sn9_79 202000.000000
Rwneg9_80 in9_80 sn9_80 78000.000000
Rwneg9_81 in9_81 sn9_81 78000.000000
Rwneg9_82 in9_82 sn9_82 202000.000000
Rwneg9_83 in9_83 sn9_83 78000.000000
Rwneg9_84 in9_84 sn9_84 202000.000000
Rwneg10_1 in10_1 sn10_1 202000.000000
Rwneg10_2 in10_2 sn10_2 78000.000000
Rwneg10_3 in10_3 sn10_3 78000.000000
Rwneg10_4 in10_4 sn10_4 202000.000000
Rwneg10_5 in10_5 sn10_5 78000.000000
Rwneg10_6 in10_6 sn10_6 202000.000000
Rwneg10_7 in10_7 sn10_7 202000.000000
Rwneg10_8 in10_8 sn10_8 78000.000000
Rwneg10_9 in10_9 sn10_9 202000.000000
Rwneg10_10 in10_10 sn10_10 78000.000000
Rwneg10_11 in10_11 sn10_11 202000.000000
Rwneg10_12 in10_12 sn10_12 78000.000000
Rwneg10_13 in10_13 sn10_13 202000.000000
Rwneg10_14 in10_14 sn10_14 202000.000000
Rwneg10_15 in10_15 sn10_15 78000.000000
Rwneg10_16 in10_16 sn10_16 202000.000000
Rwneg10_17 in10_17 sn10_17 202000.000000
Rwneg10_18 in10_18 sn10_18 78000.000000
Rwneg10_19 in10_19 sn10_19 202000.000000
Rwneg10_20 in10_20 sn10_20 202000.000000
Rwneg10_21 in10_21 sn10_21 78000.000000
Rwneg10_22 in10_22 sn10_22 78000.000000
Rwneg10_23 in10_23 sn10_23 78000.000000
Rwneg10_24 in10_24 sn10_24 78000.000000
Rwneg10_25 in10_25 sn10_25 202000.000000
Rwneg10_26 in10_26 sn10_26 78000.000000
Rwneg10_27 in10_27 sn10_27 202000.000000
Rwneg10_28 in10_28 sn10_28 202000.000000
Rwneg10_29 in10_29 sn10_29 78000.000000
Rwneg10_30 in10_30 sn10_30 202000.000000
Rwneg10_31 in10_31 sn10_31 202000.000000
Rwneg10_32 in10_32 sn10_32 78000.000000
Rwneg10_33 in10_33 sn10_33 78000.000000
Rwneg10_34 in10_34 sn10_34 202000.000000
Rwneg10_35 in10_35 sn10_35 78000.000000
Rwneg10_36 in10_36 sn10_36 78000.000000
Rwneg10_37 in10_37 sn10_37 202000.000000
Rwneg10_38 in10_38 sn10_38 202000.000000
Rwneg10_39 in10_39 sn10_39 202000.000000
Rwneg10_40 in10_40 sn10_40 202000.000000
Rwneg10_41 in10_41 sn10_41 78000.000000
Rwneg10_42 in10_42 sn10_42 78000.000000
Rwneg10_43 in10_43 sn10_43 202000.000000
Rwneg10_44 in10_44 sn10_44 78000.000000
Rwneg10_45 in10_45 sn10_45 78000.000000
Rwneg10_46 in10_46 sn10_46 202000.000000
Rwneg10_47 in10_47 sn10_47 202000.000000
Rwneg10_48 in10_48 sn10_48 202000.000000
Rwneg10_49 in10_49 sn10_49 202000.000000
Rwneg10_50 in10_50 sn10_50 202000.000000
Rwneg10_51 in10_51 sn10_51 202000.000000
Rwneg10_52 in10_52 sn10_52 202000.000000
Rwneg10_53 in10_53 sn10_53 202000.000000
Rwneg10_54 in10_54 sn10_54 202000.000000
Rwneg10_55 in10_55 sn10_55 202000.000000
Rwneg10_56 in10_56 sn10_56 78000.000000
Rwneg10_57 in10_57 sn10_57 78000.000000
Rwneg10_58 in10_58 sn10_58 78000.000000
Rwneg10_59 in10_59 sn10_59 78000.000000
Rwneg10_60 in10_60 sn10_60 78000.000000
Rwneg10_61 in10_61 sn10_61 78000.000000
Rwneg10_62 in10_62 sn10_62 202000.000000
Rwneg10_63 in10_63 sn10_63 78000.000000
Rwneg10_64 in10_64 sn10_64 202000.000000
Rwneg10_65 in10_65 sn10_65 78000.000000
Rwneg10_66 in10_66 sn10_66 78000.000000
Rwneg10_67 in10_67 sn10_67 202000.000000
Rwneg10_68 in10_68 sn10_68 202000.000000
Rwneg10_69 in10_69 sn10_69 78000.000000
Rwneg10_70 in10_70 sn10_70 78000.000000
Rwneg10_71 in10_71 sn10_71 78000.000000
Rwneg10_72 in10_72 sn10_72 78000.000000
Rwneg10_73 in10_73 sn10_73 78000.000000
Rwneg10_74 in10_74 sn10_74 202000.000000
Rwneg10_75 in10_75 sn10_75 78000.000000
Rwneg10_76 in10_76 sn10_76 78000.000000
Rwneg10_77 in10_77 sn10_77 78000.000000
Rwneg10_78 in10_78 sn10_78 78000.000000
Rwneg10_79 in10_79 sn10_79 202000.000000
Rwneg10_80 in10_80 sn10_80 78000.000000
Rwneg10_81 in10_81 sn10_81 78000.000000
Rwneg10_82 in10_82 sn10_82 78000.000000
Rwneg10_83 in10_83 sn10_83 78000.000000
Rwneg10_84 in10_84 sn10_84 78000.000000
Rwneg11_1 in11_1 sn11_1 202000.000000
Rwneg11_2 in11_2 sn11_2 202000.000000
Rwneg11_3 in11_3 sn11_3 202000.000000
Rwneg11_4 in11_4 sn11_4 202000.000000
Rwneg11_5 in11_5 sn11_5 202000.000000
Rwneg11_6 in11_6 sn11_6 78000.000000
Rwneg11_7 in11_7 sn11_7 78000.000000
Rwneg11_8 in11_8 sn11_8 202000.000000
Rwneg11_9 in11_9 sn11_9 202000.000000
Rwneg11_10 in11_10 sn11_10 78000.000000
Rwneg11_11 in11_11 sn11_11 78000.000000
Rwneg11_12 in11_12 sn11_12 202000.000000
Rwneg11_13 in11_13 sn11_13 202000.000000
Rwneg11_14 in11_14 sn11_14 78000.000000
Rwneg11_15 in11_15 sn11_15 202000.000000
Rwneg11_16 in11_16 sn11_16 202000.000000
Rwneg11_17 in11_17 sn11_17 78000.000000
Rwneg11_18 in11_18 sn11_18 202000.000000
Rwneg11_19 in11_19 sn11_19 202000.000000
Rwneg11_20 in11_20 sn11_20 202000.000000
Rwneg11_21 in11_21 sn11_21 202000.000000
Rwneg11_22 in11_22 sn11_22 202000.000000
Rwneg11_23 in11_23 sn11_23 202000.000000
Rwneg11_24 in11_24 sn11_24 78000.000000
Rwneg11_25 in11_25 sn11_25 78000.000000
Rwneg11_26 in11_26 sn11_26 202000.000000
Rwneg11_27 in11_27 sn11_27 202000.000000
Rwneg11_28 in11_28 sn11_28 202000.000000
Rwneg11_29 in11_29 sn11_29 78000.000000
Rwneg11_30 in11_30 sn11_30 202000.000000
Rwneg11_31 in11_31 sn11_31 78000.000000
Rwneg11_32 in11_32 sn11_32 202000.000000
Rwneg11_33 in11_33 sn11_33 202000.000000
Rwneg11_34 in11_34 sn11_34 78000.000000
Rwneg11_35 in11_35 sn11_35 202000.000000
Rwneg11_36 in11_36 sn11_36 78000.000000
Rwneg11_37 in11_37 sn11_37 78000.000000
Rwneg11_38 in11_38 sn11_38 202000.000000
Rwneg11_39 in11_39 sn11_39 202000.000000
Rwneg11_40 in11_40 sn11_40 202000.000000
Rwneg11_41 in11_41 sn11_41 202000.000000
Rwneg11_42 in11_42 sn11_42 202000.000000
Rwneg11_43 in11_43 sn11_43 202000.000000
Rwneg11_44 in11_44 sn11_44 78000.000000
Rwneg11_45 in11_45 sn11_45 202000.000000
Rwneg11_46 in11_46 sn11_46 78000.000000
Rwneg11_47 in11_47 sn11_47 202000.000000
Rwneg11_48 in11_48 sn11_48 78000.000000
Rwneg11_49 in11_49 sn11_49 78000.000000
Rwneg11_50 in11_50 sn11_50 78000.000000
Rwneg11_51 in11_51 sn11_51 78000.000000
Rwneg11_52 in11_52 sn11_52 202000.000000
Rwneg11_53 in11_53 sn11_53 78000.000000
Rwneg11_54 in11_54 sn11_54 202000.000000
Rwneg11_55 in11_55 sn11_55 202000.000000
Rwneg11_56 in11_56 sn11_56 78000.000000
Rwneg11_57 in11_57 sn11_57 78000.000000
Rwneg11_58 in11_58 sn11_58 202000.000000
Rwneg11_59 in11_59 sn11_59 78000.000000
Rwneg11_60 in11_60 sn11_60 78000.000000
Rwneg11_61 in11_61 sn11_61 202000.000000
Rwneg11_62 in11_62 sn11_62 78000.000000
Rwneg11_63 in11_63 sn11_63 202000.000000
Rwneg11_64 in11_64 sn11_64 78000.000000
Rwneg11_65 in11_65 sn11_65 78000.000000
Rwneg11_66 in11_66 sn11_66 78000.000000
Rwneg11_67 in11_67 sn11_67 202000.000000
Rwneg11_68 in11_68 sn11_68 202000.000000
Rwneg11_69 in11_69 sn11_69 78000.000000
Rwneg11_70 in11_70 sn11_70 78000.000000
Rwneg11_71 in11_71 sn11_71 78000.000000
Rwneg11_72 in11_72 sn11_72 202000.000000
Rwneg11_73 in11_73 sn11_73 78000.000000
Rwneg11_74 in11_74 sn11_74 202000.000000
Rwneg11_75 in11_75 sn11_75 78000.000000
Rwneg11_76 in11_76 sn11_76 202000.000000
Rwneg11_77 in11_77 sn11_77 202000.000000
Rwneg11_78 in11_78 sn11_78 202000.000000
Rwneg11_79 in11_79 sn11_79 78000.000000
Rwneg11_80 in11_80 sn11_80 202000.000000
Rwneg11_81 in11_81 sn11_81 78000.000000
Rwneg11_82 in11_82 sn11_82 202000.000000
Rwneg11_83 in11_83 sn11_83 202000.000000
Rwneg11_84 in11_84 sn11_84 202000.000000
Rwneg12_1 in12_1 sn12_1 78000.000000
Rwneg12_2 in12_2 sn12_2 78000.000000
Rwneg12_3 in12_3 sn12_3 78000.000000
Rwneg12_4 in12_4 sn12_4 202000.000000
Rwneg12_5 in12_5 sn12_5 78000.000000
Rwneg12_6 in12_6 sn12_6 202000.000000
Rwneg12_7 in12_7 sn12_7 78000.000000
Rwneg12_8 in12_8 sn12_8 202000.000000
Rwneg12_9 in12_9 sn12_9 202000.000000
Rwneg12_10 in12_10 sn12_10 202000.000000
Rwneg12_11 in12_11 sn12_11 202000.000000
Rwneg12_12 in12_12 sn12_12 202000.000000
Rwneg12_13 in12_13 sn12_13 202000.000000
Rwneg12_14 in12_14 sn12_14 78000.000000
Rwneg12_15 in12_15 sn12_15 202000.000000
Rwneg12_16 in12_16 sn12_16 202000.000000
Rwneg12_17 in12_17 sn12_17 78000.000000
Rwneg12_18 in12_18 sn12_18 202000.000000
Rwneg12_19 in12_19 sn12_19 202000.000000
Rwneg12_20 in12_20 sn12_20 202000.000000
Rwneg12_21 in12_21 sn12_21 202000.000000
Rwneg12_22 in12_22 sn12_22 202000.000000
Rwneg12_23 in12_23 sn12_23 202000.000000
Rwneg12_24 in12_24 sn12_24 78000.000000
Rwneg12_25 in12_25 sn12_25 78000.000000
Rwneg12_26 in12_26 sn12_26 78000.000000
Rwneg12_27 in12_27 sn12_27 78000.000000
Rwneg12_28 in12_28 sn12_28 78000.000000
Rwneg12_29 in12_29 sn12_29 202000.000000
Rwneg12_30 in12_30 sn12_30 202000.000000
Rwneg12_31 in12_31 sn12_31 78000.000000
Rwneg12_32 in12_32 sn12_32 78000.000000
Rwneg12_33 in12_33 sn12_33 202000.000000
Rwneg12_34 in12_34 sn12_34 202000.000000
Rwneg12_35 in12_35 sn12_35 78000.000000
Rwneg12_36 in12_36 sn12_36 78000.000000
Rwneg12_37 in12_37 sn12_37 202000.000000
Rwneg12_38 in12_38 sn12_38 202000.000000
Rwneg12_39 in12_39 sn12_39 78000.000000
Rwneg12_40 in12_40 sn12_40 202000.000000
Rwneg12_41 in12_41 sn12_41 78000.000000
Rwneg12_42 in12_42 sn12_42 78000.000000
Rwneg12_43 in12_43 sn12_43 202000.000000
Rwneg12_44 in12_44 sn12_44 78000.000000
Rwneg12_45 in12_45 sn12_45 202000.000000
Rwneg12_46 in12_46 sn12_46 78000.000000
Rwneg12_47 in12_47 sn12_47 78000.000000
Rwneg12_48 in12_48 sn12_48 78000.000000
Rwneg12_49 in12_49 sn12_49 202000.000000
Rwneg12_50 in12_50 sn12_50 78000.000000
Rwneg12_51 in12_51 sn12_51 202000.000000
Rwneg12_52 in12_52 sn12_52 202000.000000
Rwneg12_53 in12_53 sn12_53 78000.000000
Rwneg12_54 in12_54 sn12_54 78000.000000
Rwneg12_55 in12_55 sn12_55 78000.000000
Rwneg12_56 in12_56 sn12_56 202000.000000
Rwneg12_57 in12_57 sn12_57 202000.000000
Rwneg12_58 in12_58 sn12_58 202000.000000
Rwneg12_59 in12_59 sn12_59 202000.000000
Rwneg12_60 in12_60 sn12_60 78000.000000
Rwneg12_61 in12_61 sn12_61 202000.000000
Rwneg12_62 in12_62 sn12_62 78000.000000
Rwneg12_63 in12_63 sn12_63 202000.000000
Rwneg12_64 in12_64 sn12_64 202000.000000
Rwneg12_65 in12_65 sn12_65 78000.000000
Rwneg12_66 in12_66 sn12_66 202000.000000
Rwneg12_67 in12_67 sn12_67 78000.000000
Rwneg12_68 in12_68 sn12_68 202000.000000
Rwneg12_69 in12_69 sn12_69 202000.000000
Rwneg12_70 in12_70 sn12_70 202000.000000
Rwneg12_71 in12_71 sn12_71 202000.000000
Rwneg12_72 in12_72 sn12_72 78000.000000
Rwneg12_73 in12_73 sn12_73 202000.000000
Rwneg12_74 in12_74 sn12_74 78000.000000
Rwneg12_75 in12_75 sn12_75 78000.000000
Rwneg12_76 in12_76 sn12_76 78000.000000
Rwneg12_77 in12_77 sn12_77 202000.000000
Rwneg12_78 in12_78 sn12_78 202000.000000
Rwneg12_79 in12_79 sn12_79 202000.000000
Rwneg12_80 in12_80 sn12_80 202000.000000
Rwneg12_81 in12_81 sn12_81 78000.000000
Rwneg12_82 in12_82 sn12_82 202000.000000
Rwneg12_83 in12_83 sn12_83 202000.000000
Rwneg12_84 in12_84 sn12_84 202000.000000
Rwneg13_1 in13_1 sn13_1 202000.000000
Rwneg13_2 in13_2 sn13_2 202000.000000
Rwneg13_3 in13_3 sn13_3 78000.000000
Rwneg13_4 in13_4 sn13_4 202000.000000
Rwneg13_5 in13_5 sn13_5 202000.000000
Rwneg13_6 in13_6 sn13_6 78000.000000
Rwneg13_7 in13_7 sn13_7 202000.000000
Rwneg13_8 in13_8 sn13_8 202000.000000
Rwneg13_9 in13_9 sn13_9 202000.000000
Rwneg13_10 in13_10 sn13_10 78000.000000
Rwneg13_11 in13_11 sn13_11 78000.000000
Rwneg13_12 in13_12 sn13_12 202000.000000
Rwneg13_13 in13_13 sn13_13 78000.000000
Rwneg13_14 in13_14 sn13_14 78000.000000
Rwneg13_15 in13_15 sn13_15 78000.000000
Rwneg13_16 in13_16 sn13_16 202000.000000
Rwneg13_17 in13_17 sn13_17 78000.000000
Rwneg13_18 in13_18 sn13_18 202000.000000
Rwneg13_19 in13_19 sn13_19 78000.000000
Rwneg13_20 in13_20 sn13_20 78000.000000
Rwneg13_21 in13_21 sn13_21 202000.000000
Rwneg13_22 in13_22 sn13_22 202000.000000
Rwneg13_23 in13_23 sn13_23 78000.000000
Rwneg13_24 in13_24 sn13_24 78000.000000
Rwneg13_25 in13_25 sn13_25 202000.000000
Rwneg13_26 in13_26 sn13_26 78000.000000
Rwneg13_27 in13_27 sn13_27 202000.000000
Rwneg13_28 in13_28 sn13_28 78000.000000
Rwneg13_29 in13_29 sn13_29 202000.000000
Rwneg13_30 in13_30 sn13_30 202000.000000
Rwneg13_31 in13_31 sn13_31 202000.000000
Rwneg13_32 in13_32 sn13_32 78000.000000
Rwneg13_33 in13_33 sn13_33 78000.000000
Rwneg13_34 in13_34 sn13_34 78000.000000
Rwneg13_35 in13_35 sn13_35 202000.000000
Rwneg13_36 in13_36 sn13_36 202000.000000
Rwneg13_37 in13_37 sn13_37 202000.000000
Rwneg13_38 in13_38 sn13_38 78000.000000
Rwneg13_39 in13_39 sn13_39 78000.000000
Rwneg13_40 in13_40 sn13_40 78000.000000
Rwneg13_41 in13_41 sn13_41 202000.000000
Rwneg13_42 in13_42 sn13_42 202000.000000
Rwneg13_43 in13_43 sn13_43 202000.000000
Rwneg13_44 in13_44 sn13_44 202000.000000
Rwneg13_45 in13_45 sn13_45 78000.000000
Rwneg13_46 in13_46 sn13_46 78000.000000
Rwneg13_47 in13_47 sn13_47 78000.000000
Rwneg13_48 in13_48 sn13_48 78000.000000
Rwneg13_49 in13_49 sn13_49 202000.000000
Rwneg13_50 in13_50 sn13_50 78000.000000
Rwneg13_51 in13_51 sn13_51 202000.000000
Rwneg13_52 in13_52 sn13_52 202000.000000
Rwneg13_53 in13_53 sn13_53 202000.000000
Rwneg13_54 in13_54 sn13_54 202000.000000
Rwneg13_55 in13_55 sn13_55 78000.000000
Rwneg13_56 in13_56 sn13_56 202000.000000
Rwneg13_57 in13_57 sn13_57 202000.000000
Rwneg13_58 in13_58 sn13_58 78000.000000
Rwneg13_59 in13_59 sn13_59 202000.000000
Rwneg13_60 in13_60 sn13_60 202000.000000
Rwneg13_61 in13_61 sn13_61 202000.000000
Rwneg13_62 in13_62 sn13_62 202000.000000
Rwneg13_63 in13_63 sn13_63 202000.000000
Rwneg13_64 in13_64 sn13_64 202000.000000
Rwneg13_65 in13_65 sn13_65 202000.000000
Rwneg13_66 in13_66 sn13_66 202000.000000
Rwneg13_67 in13_67 sn13_67 78000.000000
Rwneg13_68 in13_68 sn13_68 202000.000000
Rwneg13_69 in13_69 sn13_69 202000.000000
Rwneg13_70 in13_70 sn13_70 202000.000000
Rwneg13_71 in13_71 sn13_71 202000.000000
Rwneg13_72 in13_72 sn13_72 202000.000000
Rwneg13_73 in13_73 sn13_73 202000.000000
Rwneg13_74 in13_74 sn13_74 78000.000000
Rwneg13_75 in13_75 sn13_75 78000.000000
Rwneg13_76 in13_76 sn13_76 202000.000000
Rwneg13_77 in13_77 sn13_77 78000.000000
Rwneg13_78 in13_78 sn13_78 202000.000000
Rwneg13_79 in13_79 sn13_79 202000.000000
Rwneg13_80 in13_80 sn13_80 202000.000000
Rwneg13_81 in13_81 sn13_81 78000.000000
Rwneg13_82 in13_82 sn13_82 202000.000000
Rwneg13_83 in13_83 sn13_83 78000.000000
Rwneg13_84 in13_84 sn13_84 202000.000000
Rwneg14_1 in14_1 sn14_1 202000.000000
Rwneg14_2 in14_2 sn14_2 202000.000000
Rwneg14_3 in14_3 sn14_3 202000.000000
Rwneg14_4 in14_4 sn14_4 78000.000000
Rwneg14_5 in14_5 sn14_5 78000.000000
Rwneg14_6 in14_6 sn14_6 202000.000000
Rwneg14_7 in14_7 sn14_7 202000.000000
Rwneg14_8 in14_8 sn14_8 78000.000000
Rwneg14_9 in14_9 sn14_9 78000.000000
Rwneg14_10 in14_10 sn14_10 78000.000000
Rwneg14_11 in14_11 sn14_11 202000.000000
Rwneg14_12 in14_12 sn14_12 78000.000000
Rwneg14_13 in14_13 sn14_13 78000.000000
Rwneg14_14 in14_14 sn14_14 202000.000000
Rwneg14_15 in14_15 sn14_15 78000.000000
Rwneg14_16 in14_16 sn14_16 202000.000000
Rwneg14_17 in14_17 sn14_17 202000.000000
Rwneg14_18 in14_18 sn14_18 78000.000000
Rwneg14_19 in14_19 sn14_19 202000.000000
Rwneg14_20 in14_20 sn14_20 78000.000000
Rwneg14_21 in14_21 sn14_21 202000.000000
Rwneg14_22 in14_22 sn14_22 202000.000000
Rwneg14_23 in14_23 sn14_23 202000.000000
Rwneg14_24 in14_24 sn14_24 78000.000000
Rwneg14_25 in14_25 sn14_25 202000.000000
Rwneg14_26 in14_26 sn14_26 202000.000000
Rwneg14_27 in14_27 sn14_27 78000.000000
Rwneg14_28 in14_28 sn14_28 78000.000000
Rwneg14_29 in14_29 sn14_29 202000.000000
Rwneg14_30 in14_30 sn14_30 202000.000000
Rwneg14_31 in14_31 sn14_31 202000.000000
Rwneg14_32 in14_32 sn14_32 78000.000000
Rwneg14_33 in14_33 sn14_33 202000.000000
Rwneg14_34 in14_34 sn14_34 202000.000000
Rwneg14_35 in14_35 sn14_35 78000.000000
Rwneg14_36 in14_36 sn14_36 78000.000000
Rwneg14_37 in14_37 sn14_37 202000.000000
Rwneg14_38 in14_38 sn14_38 202000.000000
Rwneg14_39 in14_39 sn14_39 78000.000000
Rwneg14_40 in14_40 sn14_40 202000.000000
Rwneg14_41 in14_41 sn14_41 78000.000000
Rwneg14_42 in14_42 sn14_42 202000.000000
Rwneg14_43 in14_43 sn14_43 202000.000000
Rwneg14_44 in14_44 sn14_44 202000.000000
Rwneg14_45 in14_45 sn14_45 78000.000000
Rwneg14_46 in14_46 sn14_46 202000.000000
Rwneg14_47 in14_47 sn14_47 202000.000000
Rwneg14_48 in14_48 sn14_48 78000.000000
Rwneg14_49 in14_49 sn14_49 202000.000000
Rwneg14_50 in14_50 sn14_50 202000.000000
Rwneg14_51 in14_51 sn14_51 202000.000000
Rwneg14_52 in14_52 sn14_52 202000.000000
Rwneg14_53 in14_53 sn14_53 202000.000000
Rwneg14_54 in14_54 sn14_54 78000.000000
Rwneg14_55 in14_55 sn14_55 202000.000000
Rwneg14_56 in14_56 sn14_56 78000.000000
Rwneg14_57 in14_57 sn14_57 202000.000000
Rwneg14_58 in14_58 sn14_58 202000.000000
Rwneg14_59 in14_59 sn14_59 202000.000000
Rwneg14_60 in14_60 sn14_60 78000.000000
Rwneg14_61 in14_61 sn14_61 202000.000000
Rwneg14_62 in14_62 sn14_62 202000.000000
Rwneg14_63 in14_63 sn14_63 78000.000000
Rwneg14_64 in14_64 sn14_64 202000.000000
Rwneg14_65 in14_65 sn14_65 78000.000000
Rwneg14_66 in14_66 sn14_66 202000.000000
Rwneg14_67 in14_67 sn14_67 78000.000000
Rwneg14_68 in14_68 sn14_68 78000.000000
Rwneg14_69 in14_69 sn14_69 78000.000000
Rwneg14_70 in14_70 sn14_70 78000.000000
Rwneg14_71 in14_71 sn14_71 78000.000000
Rwneg14_72 in14_72 sn14_72 202000.000000
Rwneg14_73 in14_73 sn14_73 202000.000000
Rwneg14_74 in14_74 sn14_74 202000.000000
Rwneg14_75 in14_75 sn14_75 78000.000000
Rwneg14_76 in14_76 sn14_76 202000.000000
Rwneg14_77 in14_77 sn14_77 202000.000000
Rwneg14_78 in14_78 sn14_78 202000.000000
Rwneg14_79 in14_79 sn14_79 78000.000000
Rwneg14_80 in14_80 sn14_80 78000.000000
Rwneg14_81 in14_81 sn14_81 78000.000000
Rwneg14_82 in14_82 sn14_82 78000.000000
Rwneg14_83 in14_83 sn14_83 202000.000000
Rwneg14_84 in14_84 sn14_84 78000.000000
Rwneg15_1 in15_1 sn15_1 202000.000000
Rwneg15_2 in15_2 sn15_2 202000.000000
Rwneg15_3 in15_3 sn15_3 202000.000000
Rwneg15_4 in15_4 sn15_4 78000.000000
Rwneg15_5 in15_5 sn15_5 78000.000000
Rwneg15_6 in15_6 sn15_6 202000.000000
Rwneg15_7 in15_7 sn15_7 202000.000000
Rwneg15_8 in15_8 sn15_8 78000.000000
Rwneg15_9 in15_9 sn15_9 78000.000000
Rwneg15_10 in15_10 sn15_10 78000.000000
Rwneg15_11 in15_11 sn15_11 202000.000000
Rwneg15_12 in15_12 sn15_12 202000.000000
Rwneg15_13 in15_13 sn15_13 78000.000000
Rwneg15_14 in15_14 sn15_14 78000.000000
Rwneg15_15 in15_15 sn15_15 202000.000000
Rwneg15_16 in15_16 sn15_16 202000.000000
Rwneg15_17 in15_17 sn15_17 202000.000000
Rwneg15_18 in15_18 sn15_18 78000.000000
Rwneg15_19 in15_19 sn15_19 202000.000000
Rwneg15_20 in15_20 sn15_20 78000.000000
Rwneg15_21 in15_21 sn15_21 202000.000000
Rwneg15_22 in15_22 sn15_22 202000.000000
Rwneg15_23 in15_23 sn15_23 78000.000000
Rwneg15_24 in15_24 sn15_24 202000.000000
Rwneg15_25 in15_25 sn15_25 202000.000000
Rwneg15_26 in15_26 sn15_26 78000.000000
Rwneg15_27 in15_27 sn15_27 78000.000000
Rwneg15_28 in15_28 sn15_28 202000.000000
Rwneg15_29 in15_29 sn15_29 202000.000000
Rwneg15_30 in15_30 sn15_30 78000.000000
Rwneg15_31 in15_31 sn15_31 78000.000000
Rwneg15_32 in15_32 sn15_32 78000.000000
Rwneg15_33 in15_33 sn15_33 202000.000000
Rwneg15_34 in15_34 sn15_34 202000.000000
Rwneg15_35 in15_35 sn15_35 202000.000000
Rwneg15_36 in15_36 sn15_36 202000.000000
Rwneg15_37 in15_37 sn15_37 202000.000000
Rwneg15_38 in15_38 sn15_38 78000.000000
Rwneg15_39 in15_39 sn15_39 78000.000000
Rwneg15_40 in15_40 sn15_40 202000.000000
Rwneg15_41 in15_41 sn15_41 78000.000000
Rwneg15_42 in15_42 sn15_42 202000.000000
Rwneg15_43 in15_43 sn15_43 202000.000000
Rwneg15_44 in15_44 sn15_44 202000.000000
Rwneg15_45 in15_45 sn15_45 202000.000000
Rwneg15_46 in15_46 sn15_46 78000.000000
Rwneg15_47 in15_47 sn15_47 202000.000000
Rwneg15_48 in15_48 sn15_48 78000.000000
Rwneg15_49 in15_49 sn15_49 202000.000000
Rwneg15_50 in15_50 sn15_50 78000.000000
Rwneg15_51 in15_51 sn15_51 202000.000000
Rwneg15_52 in15_52 sn15_52 202000.000000
Rwneg15_53 in15_53 sn15_53 78000.000000
Rwneg15_54 in15_54 sn15_54 78000.000000
Rwneg15_55 in15_55 sn15_55 78000.000000
Rwneg15_56 in15_56 sn15_56 202000.000000
Rwneg15_57 in15_57 sn15_57 202000.000000
Rwneg15_58 in15_58 sn15_58 202000.000000
Rwneg15_59 in15_59 sn15_59 78000.000000
Rwneg15_60 in15_60 sn15_60 202000.000000
Rwneg15_61 in15_61 sn15_61 202000.000000
Rwneg15_62 in15_62 sn15_62 78000.000000
Rwneg15_63 in15_63 sn15_63 202000.000000
Rwneg15_64 in15_64 sn15_64 78000.000000
Rwneg15_65 in15_65 sn15_65 78000.000000
Rwneg15_66 in15_66 sn15_66 202000.000000
Rwneg15_67 in15_67 sn15_67 202000.000000
Rwneg15_68 in15_68 sn15_68 202000.000000
Rwneg15_69 in15_69 sn15_69 202000.000000
Rwneg15_70 in15_70 sn15_70 202000.000000
Rwneg15_71 in15_71 sn15_71 202000.000000
Rwneg15_72 in15_72 sn15_72 202000.000000
Rwneg15_73 in15_73 sn15_73 202000.000000
Rwneg15_74 in15_74 sn15_74 202000.000000
Rwneg15_75 in15_75 sn15_75 202000.000000
Rwneg15_76 in15_76 sn15_76 202000.000000
Rwneg15_77 in15_77 sn15_77 78000.000000
Rwneg15_78 in15_78 sn15_78 202000.000000
Rwneg15_79 in15_79 sn15_79 202000.000000
Rwneg15_80 in15_80 sn15_80 78000.000000
Rwneg15_81 in15_81 sn15_81 202000.000000
Rwneg15_82 in15_82 sn15_82 78000.000000
Rwneg15_83 in15_83 sn15_83 202000.000000
Rwneg15_84 in15_84 sn15_84 78000.000000
Rwneg16_1 in16_1 sn16_1 78000.000000
Rwneg16_2 in16_2 sn16_2 78000.000000
Rwneg16_3 in16_3 sn16_3 78000.000000
Rwneg16_4 in16_4 sn16_4 202000.000000
Rwneg16_5 in16_5 sn16_5 202000.000000
Rwneg16_6 in16_6 sn16_6 202000.000000
Rwneg16_7 in16_7 sn16_7 202000.000000
Rwneg16_8 in16_8 sn16_8 78000.000000
Rwneg16_9 in16_9 sn16_9 78000.000000
Rwneg16_10 in16_10 sn16_10 202000.000000
Rwneg16_11 in16_11 sn16_11 202000.000000
Rwneg16_12 in16_12 sn16_12 202000.000000
Rwneg16_13 in16_13 sn16_13 78000.000000
Rwneg16_14 in16_14 sn16_14 202000.000000
Rwneg16_15 in16_15 sn16_15 202000.000000
Rwneg16_16 in16_16 sn16_16 202000.000000
Rwneg16_17 in16_17 sn16_17 202000.000000
Rwneg16_18 in16_18 sn16_18 78000.000000
Rwneg16_19 in16_19 sn16_19 202000.000000
Rwneg16_20 in16_20 sn16_20 202000.000000
Rwneg16_21 in16_21 sn16_21 202000.000000
Rwneg16_22 in16_22 sn16_22 202000.000000
Rwneg16_23 in16_23 sn16_23 202000.000000
Rwneg16_24 in16_24 sn16_24 78000.000000
Rwneg16_25 in16_25 sn16_25 202000.000000
Rwneg16_26 in16_26 sn16_26 78000.000000
Rwneg16_27 in16_27 sn16_27 202000.000000
Rwneg16_28 in16_28 sn16_28 202000.000000
Rwneg16_29 in16_29 sn16_29 78000.000000
Rwneg16_30 in16_30 sn16_30 202000.000000
Rwneg16_31 in16_31 sn16_31 202000.000000
Rwneg16_32 in16_32 sn16_32 202000.000000
Rwneg16_33 in16_33 sn16_33 78000.000000
Rwneg16_34 in16_34 sn16_34 202000.000000
Rwneg16_35 in16_35 sn16_35 78000.000000
Rwneg16_36 in16_36 sn16_36 78000.000000
Rwneg16_37 in16_37 sn16_37 202000.000000
Rwneg16_38 in16_38 sn16_38 202000.000000
Rwneg16_39 in16_39 sn16_39 78000.000000
Rwneg16_40 in16_40 sn16_40 202000.000000
Rwneg16_41 in16_41 sn16_41 202000.000000
Rwneg16_42 in16_42 sn16_42 78000.000000
Rwneg16_43 in16_43 sn16_43 202000.000000
Rwneg16_44 in16_44 sn16_44 202000.000000
Rwneg16_45 in16_45 sn16_45 202000.000000
Rwneg16_46 in16_46 sn16_46 202000.000000
Rwneg16_47 in16_47 sn16_47 78000.000000
Rwneg16_48 in16_48 sn16_48 202000.000000
Rwneg16_49 in16_49 sn16_49 78000.000000
Rwneg16_50 in16_50 sn16_50 202000.000000
Rwneg16_51 in16_51 sn16_51 202000.000000
Rwneg16_52 in16_52 sn16_52 78000.000000
Rwneg16_53 in16_53 sn16_53 78000.000000
Rwneg16_54 in16_54 sn16_54 202000.000000
Rwneg16_55 in16_55 sn16_55 78000.000000
Rwneg16_56 in16_56 sn16_56 202000.000000
Rwneg16_57 in16_57 sn16_57 202000.000000
Rwneg16_58 in16_58 sn16_58 202000.000000
Rwneg16_59 in16_59 sn16_59 202000.000000
Rwneg16_60 in16_60 sn16_60 78000.000000
Rwneg16_61 in16_61 sn16_61 78000.000000
Rwneg16_62 in16_62 sn16_62 202000.000000
Rwneg16_63 in16_63 sn16_63 78000.000000
Rwneg16_64 in16_64 sn16_64 78000.000000
Rwneg16_65 in16_65 sn16_65 202000.000000
Rwneg16_66 in16_66 sn16_66 78000.000000
Rwneg16_67 in16_67 sn16_67 78000.000000
Rwneg16_68 in16_68 sn16_68 202000.000000
Rwneg16_69 in16_69 sn16_69 202000.000000
Rwneg16_70 in16_70 sn16_70 202000.000000
Rwneg16_71 in16_71 sn16_71 202000.000000
Rwneg16_72 in16_72 sn16_72 202000.000000
Rwneg16_73 in16_73 sn16_73 202000.000000
Rwneg16_74 in16_74 sn16_74 78000.000000
Rwneg16_75 in16_75 sn16_75 202000.000000
Rwneg16_76 in16_76 sn16_76 78000.000000
Rwneg16_77 in16_77 sn16_77 202000.000000
Rwneg16_78 in16_78 sn16_78 202000.000000
Rwneg16_79 in16_79 sn16_79 202000.000000
Rwneg16_80 in16_80 sn16_80 78000.000000
Rwneg16_81 in16_81 sn16_81 202000.000000
Rwneg16_82 in16_82 sn16_82 78000.000000
Rwneg16_83 in16_83 sn16_83 78000.000000
Rwneg16_84 in16_84 sn16_84 202000.000000
Rwneg17_1 in17_1 sn17_1 202000.000000
Rwneg17_2 in17_2 sn17_2 202000.000000
Rwneg17_3 in17_3 sn17_3 78000.000000
Rwneg17_4 in17_4 sn17_4 202000.000000
Rwneg17_5 in17_5 sn17_5 202000.000000
Rwneg17_6 in17_6 sn17_6 202000.000000
Rwneg17_7 in17_7 sn17_7 78000.000000
Rwneg17_8 in17_8 sn17_8 202000.000000
Rwneg17_9 in17_9 sn17_9 202000.000000
Rwneg17_10 in17_10 sn17_10 202000.000000
Rwneg17_11 in17_11 sn17_11 78000.000000
Rwneg17_12 in17_12 sn17_12 202000.000000
Rwneg17_13 in17_13 sn17_13 202000.000000
Rwneg17_14 in17_14 sn17_14 78000.000000
Rwneg17_15 in17_15 sn17_15 78000.000000
Rwneg17_16 in17_16 sn17_16 202000.000000
Rwneg17_17 in17_17 sn17_17 78000.000000
Rwneg17_18 in17_18 sn17_18 202000.000000
Rwneg17_19 in17_19 sn17_19 202000.000000
Rwneg17_20 in17_20 sn17_20 202000.000000
Rwneg17_21 in17_21 sn17_21 202000.000000
Rwneg17_22 in17_22 sn17_22 202000.000000
Rwneg17_23 in17_23 sn17_23 202000.000000
Rwneg17_24 in17_24 sn17_24 78000.000000
Rwneg17_25 in17_25 sn17_25 78000.000000
Rwneg17_26 in17_26 sn17_26 202000.000000
Rwneg17_27 in17_27 sn17_27 202000.000000
Rwneg17_28 in17_28 sn17_28 202000.000000
Rwneg17_29 in17_29 sn17_29 202000.000000
Rwneg17_30 in17_30 sn17_30 78000.000000
Rwneg17_31 in17_31 sn17_31 78000.000000
Rwneg17_32 in17_32 sn17_32 202000.000000
Rwneg17_33 in17_33 sn17_33 78000.000000
Rwneg17_34 in17_34 sn17_34 202000.000000
Rwneg17_35 in17_35 sn17_35 78000.000000
Rwneg17_36 in17_36 sn17_36 202000.000000
Rwneg17_37 in17_37 sn17_37 202000.000000
Rwneg17_38 in17_38 sn17_38 202000.000000
Rwneg17_39 in17_39 sn17_39 202000.000000
Rwneg17_40 in17_40 sn17_40 202000.000000
Rwneg17_41 in17_41 sn17_41 202000.000000
Rwneg17_42 in17_42 sn17_42 202000.000000
Rwneg17_43 in17_43 sn17_43 78000.000000
Rwneg17_44 in17_44 sn17_44 202000.000000
Rwneg17_45 in17_45 sn17_45 202000.000000
Rwneg17_46 in17_46 sn17_46 78000.000000
Rwneg17_47 in17_47 sn17_47 78000.000000
Rwneg17_48 in17_48 sn17_48 202000.000000
Rwneg17_49 in17_49 sn17_49 78000.000000
Rwneg17_50 in17_50 sn17_50 78000.000000
Rwneg17_51 in17_51 sn17_51 78000.000000
Rwneg17_52 in17_52 sn17_52 78000.000000
Rwneg17_53 in17_53 sn17_53 78000.000000
Rwneg17_54 in17_54 sn17_54 78000.000000
Rwneg17_55 in17_55 sn17_55 202000.000000
Rwneg17_56 in17_56 sn17_56 202000.000000
Rwneg17_57 in17_57 sn17_57 78000.000000
Rwneg17_58 in17_58 sn17_58 202000.000000
Rwneg17_59 in17_59 sn17_59 78000.000000
Rwneg17_60 in17_60 sn17_60 202000.000000
Rwneg17_61 in17_61 sn17_61 202000.000000
Rwneg17_62 in17_62 sn17_62 78000.000000
Rwneg17_63 in17_63 sn17_63 202000.000000
Rwneg17_64 in17_64 sn17_64 202000.000000
Rwneg17_65 in17_65 sn17_65 202000.000000
Rwneg17_66 in17_66 sn17_66 202000.000000
Rwneg17_67 in17_67 sn17_67 78000.000000
Rwneg17_68 in17_68 sn17_68 202000.000000
Rwneg17_69 in17_69 sn17_69 78000.000000
Rwneg17_70 in17_70 sn17_70 202000.000000
Rwneg17_71 in17_71 sn17_71 202000.000000
Rwneg17_72 in17_72 sn17_72 78000.000000
Rwneg17_73 in17_73 sn17_73 202000.000000
Rwneg17_74 in17_74 sn17_74 78000.000000
Rwneg17_75 in17_75 sn17_75 78000.000000
Rwneg17_76 in17_76 sn17_76 78000.000000
Rwneg17_77 in17_77 sn17_77 202000.000000
Rwneg17_78 in17_78 sn17_78 202000.000000
Rwneg17_79 in17_79 sn17_79 202000.000000
Rwneg17_80 in17_80 sn17_80 202000.000000
Rwneg17_81 in17_81 sn17_81 78000.000000
Rwneg17_82 in17_82 sn17_82 202000.000000
Rwneg17_83 in17_83 sn17_83 202000.000000
Rwneg17_84 in17_84 sn17_84 202000.000000
Rwneg18_1 in18_1 sn18_1 78000.000000
Rwneg18_2 in18_2 sn18_2 202000.000000
Rwneg18_3 in18_3 sn18_3 202000.000000
Rwneg18_4 in18_4 sn18_4 78000.000000
Rwneg18_5 in18_5 sn18_5 78000.000000
Rwneg18_6 in18_6 sn18_6 78000.000000
Rwneg18_7 in18_7 sn18_7 202000.000000
Rwneg18_8 in18_8 sn18_8 202000.000000
Rwneg18_9 in18_9 sn18_9 78000.000000
Rwneg18_10 in18_10 sn18_10 202000.000000
Rwneg18_11 in18_11 sn18_11 202000.000000
Rwneg18_12 in18_12 sn18_12 78000.000000
Rwneg18_13 in18_13 sn18_13 78000.000000
Rwneg18_14 in18_14 sn18_14 78000.000000
Rwneg18_15 in18_15 sn18_15 78000.000000
Rwneg18_16 in18_16 sn18_16 78000.000000
Rwneg18_17 in18_17 sn18_17 78000.000000
Rwneg18_18 in18_18 sn18_18 78000.000000
Rwneg18_19 in18_19 sn18_19 78000.000000
Rwneg18_20 in18_20 sn18_20 78000.000000
Rwneg18_21 in18_21 sn18_21 202000.000000
Rwneg18_22 in18_22 sn18_22 78000.000000
Rwneg18_23 in18_23 sn18_23 202000.000000
Rwneg18_24 in18_24 sn18_24 78000.000000
Rwneg18_25 in18_25 sn18_25 202000.000000
Rwneg18_26 in18_26 sn18_26 78000.000000
Rwneg18_27 in18_27 sn18_27 78000.000000
Rwneg18_28 in18_28 sn18_28 78000.000000
Rwneg18_29 in18_29 sn18_29 78000.000000
Rwneg18_30 in18_30 sn18_30 78000.000000
Rwneg18_31 in18_31 sn18_31 78000.000000
Rwneg18_32 in18_32 sn18_32 78000.000000
Rwneg18_33 in18_33 sn18_33 202000.000000
Rwneg18_34 in18_34 sn18_34 78000.000000
Rwneg18_35 in18_35 sn18_35 78000.000000
Rwneg18_36 in18_36 sn18_36 78000.000000
Rwneg18_37 in18_37 sn18_37 202000.000000
Rwneg18_38 in18_38 sn18_38 78000.000000
Rwneg18_39 in18_39 sn18_39 78000.000000
Rwneg18_40 in18_40 sn18_40 202000.000000
Rwneg18_41 in18_41 sn18_41 202000.000000
Rwneg18_42 in18_42 sn18_42 202000.000000
Rwneg18_43 in18_43 sn18_43 202000.000000
Rwneg18_44 in18_44 sn18_44 202000.000000
Rwneg18_45 in18_45 sn18_45 78000.000000
Rwneg18_46 in18_46 sn18_46 202000.000000
Rwneg18_47 in18_47 sn18_47 78000.000000
Rwneg18_48 in18_48 sn18_48 78000.000000
Rwneg18_49 in18_49 sn18_49 202000.000000
Rwneg18_50 in18_50 sn18_50 202000.000000
Rwneg18_51 in18_51 sn18_51 202000.000000
Rwneg18_52 in18_52 sn18_52 202000.000000
Rwneg18_53 in18_53 sn18_53 202000.000000
Rwneg18_54 in18_54 sn18_54 78000.000000
Rwneg18_55 in18_55 sn18_55 78000.000000
Rwneg18_56 in18_56 sn18_56 78000.000000
Rwneg18_57 in18_57 sn18_57 78000.000000
Rwneg18_58 in18_58 sn18_58 202000.000000
Rwneg18_59 in18_59 sn18_59 78000.000000
Rwneg18_60 in18_60 sn18_60 202000.000000
Rwneg18_61 in18_61 sn18_61 202000.000000
Rwneg18_62 in18_62 sn18_62 78000.000000
Rwneg18_63 in18_63 sn18_63 202000.000000
Rwneg18_64 in18_64 sn18_64 78000.000000
Rwneg18_65 in18_65 sn18_65 78000.000000
Rwneg18_66 in18_66 sn18_66 202000.000000
Rwneg18_67 in18_67 sn18_67 78000.000000
Rwneg18_68 in18_68 sn18_68 78000.000000
Rwneg18_69 in18_69 sn18_69 78000.000000
Rwneg18_70 in18_70 sn18_70 202000.000000
Rwneg18_71 in18_71 sn18_71 78000.000000
Rwneg18_72 in18_72 sn18_72 78000.000000
Rwneg18_73 in18_73 sn18_73 202000.000000
Rwneg18_74 in18_74 sn18_74 202000.000000
Rwneg18_75 in18_75 sn18_75 78000.000000
Rwneg18_76 in18_76 sn18_76 202000.000000
Rwneg18_77 in18_77 sn18_77 78000.000000
Rwneg18_78 in18_78 sn18_78 202000.000000
Rwneg18_79 in18_79 sn18_79 202000.000000
Rwneg18_80 in18_80 sn18_80 78000.000000
Rwneg18_81 in18_81 sn18_81 202000.000000
Rwneg18_82 in18_82 sn18_82 78000.000000
Rwneg18_83 in18_83 sn18_83 202000.000000
Rwneg18_84 in18_84 sn18_84 202000.000000
Rwneg19_1 in19_1 sn19_1 202000.000000
Rwneg19_2 in19_2 sn19_2 202000.000000
Rwneg19_3 in19_3 sn19_3 202000.000000
Rwneg19_4 in19_4 sn19_4 202000.000000
Rwneg19_5 in19_5 sn19_5 78000.000000
Rwneg19_6 in19_6 sn19_6 78000.000000
Rwneg19_7 in19_7 sn19_7 78000.000000
Rwneg19_8 in19_8 sn19_8 202000.000000
Rwneg19_9 in19_9 sn19_9 202000.000000
Rwneg19_10 in19_10 sn19_10 202000.000000
Rwneg19_11 in19_11 sn19_11 202000.000000
Rwneg19_12 in19_12 sn19_12 78000.000000
Rwneg19_13 in19_13 sn19_13 202000.000000
Rwneg19_14 in19_14 sn19_14 202000.000000
Rwneg19_15 in19_15 sn19_15 202000.000000
Rwneg19_16 in19_16 sn19_16 78000.000000
Rwneg19_17 in19_17 sn19_17 78000.000000
Rwneg19_18 in19_18 sn19_18 202000.000000
Rwneg19_19 in19_19 sn19_19 78000.000000
Rwneg19_20 in19_20 sn19_20 202000.000000
Rwneg19_21 in19_21 sn19_21 78000.000000
Rwneg19_22 in19_22 sn19_22 202000.000000
Rwneg19_23 in19_23 sn19_23 78000.000000
Rwneg19_24 in19_24 sn19_24 78000.000000
Rwneg19_25 in19_25 sn19_25 202000.000000
Rwneg19_26 in19_26 sn19_26 202000.000000
Rwneg19_27 in19_27 sn19_27 202000.000000
Rwneg19_28 in19_28 sn19_28 78000.000000
Rwneg19_29 in19_29 sn19_29 202000.000000
Rwneg19_30 in19_30 sn19_30 78000.000000
Rwneg19_31 in19_31 sn19_31 78000.000000
Rwneg19_32 in19_32 sn19_32 78000.000000
Rwneg19_33 in19_33 sn19_33 202000.000000
Rwneg19_34 in19_34 sn19_34 78000.000000
Rwneg19_35 in19_35 sn19_35 202000.000000
Rwneg19_36 in19_36 sn19_36 202000.000000
Rwneg19_37 in19_37 sn19_37 78000.000000
Rwneg19_38 in19_38 sn19_38 78000.000000
Rwneg19_39 in19_39 sn19_39 202000.000000
Rwneg19_40 in19_40 sn19_40 78000.000000
Rwneg19_41 in19_41 sn19_41 78000.000000
Rwneg19_42 in19_42 sn19_42 202000.000000
Rwneg19_43 in19_43 sn19_43 202000.000000
Rwneg19_44 in19_44 sn19_44 78000.000000
Rwneg19_45 in19_45 sn19_45 202000.000000
Rwneg19_46 in19_46 sn19_46 202000.000000
Rwneg19_47 in19_47 sn19_47 78000.000000
Rwneg19_48 in19_48 sn19_48 78000.000000
Rwneg19_49 in19_49 sn19_49 202000.000000
Rwneg19_50 in19_50 sn19_50 78000.000000
Rwneg19_51 in19_51 sn19_51 78000.000000
Rwneg19_52 in19_52 sn19_52 78000.000000
Rwneg19_53 in19_53 sn19_53 78000.000000
Rwneg19_54 in19_54 sn19_54 78000.000000
Rwneg19_55 in19_55 sn19_55 78000.000000
Rwneg19_56 in19_56 sn19_56 202000.000000
Rwneg19_57 in19_57 sn19_57 202000.000000
Rwneg19_58 in19_58 sn19_58 78000.000000
Rwneg19_59 in19_59 sn19_59 202000.000000
Rwneg19_60 in19_60 sn19_60 202000.000000
Rwneg19_61 in19_61 sn19_61 202000.000000
Rwneg19_62 in19_62 sn19_62 78000.000000
Rwneg19_63 in19_63 sn19_63 202000.000000
Rwneg19_64 in19_64 sn19_64 202000.000000
Rwneg19_65 in19_65 sn19_65 202000.000000
Rwneg19_66 in19_66 sn19_66 202000.000000
Rwneg19_67 in19_67 sn19_67 78000.000000
Rwneg19_68 in19_68 sn19_68 78000.000000
Rwneg19_69 in19_69 sn19_69 202000.000000
Rwneg19_70 in19_70 sn19_70 202000.000000
Rwneg19_71 in19_71 sn19_71 202000.000000
Rwneg19_72 in19_72 sn19_72 78000.000000
Rwneg19_73 in19_73 sn19_73 78000.000000
Rwneg19_74 in19_74 sn19_74 202000.000000
Rwneg19_75 in19_75 sn19_75 202000.000000
Rwneg19_76 in19_76 sn19_76 202000.000000
Rwneg19_77 in19_77 sn19_77 202000.000000
Rwneg19_78 in19_78 sn19_78 78000.000000
Rwneg19_79 in19_79 sn19_79 202000.000000
Rwneg19_80 in19_80 sn19_80 78000.000000
Rwneg19_81 in19_81 sn19_81 202000.000000
Rwneg19_82 in19_82 sn19_82 202000.000000
Rwneg19_83 in19_83 sn19_83 202000.000000
Rwneg19_84 in19_84 sn19_84 202000.000000
Rwneg20_1 in20_1 sn20_1 78000.000000
Rwneg20_2 in20_2 sn20_2 78000.000000
Rwneg20_3 in20_3 sn20_3 202000.000000
Rwneg20_4 in20_4 sn20_4 78000.000000
Rwneg20_5 in20_5 sn20_5 202000.000000
Rwneg20_6 in20_6 sn20_6 202000.000000
Rwneg20_7 in20_7 sn20_7 78000.000000
Rwneg20_8 in20_8 sn20_8 78000.000000
Rwneg20_9 in20_9 sn20_9 78000.000000
Rwneg20_10 in20_10 sn20_10 202000.000000
Rwneg20_11 in20_11 sn20_11 78000.000000
Rwneg20_12 in20_12 sn20_12 202000.000000
Rwneg20_13 in20_13 sn20_13 202000.000000
Rwneg20_14 in20_14 sn20_14 202000.000000
Rwneg20_15 in20_15 sn20_15 78000.000000
Rwneg20_16 in20_16 sn20_16 202000.000000
Rwneg20_17 in20_17 sn20_17 78000.000000
Rwneg20_18 in20_18 sn20_18 202000.000000
Rwneg20_19 in20_19 sn20_19 78000.000000
Rwneg20_20 in20_20 sn20_20 202000.000000
Rwneg20_21 in20_21 sn20_21 78000.000000
Rwneg20_22 in20_22 sn20_22 202000.000000
Rwneg20_23 in20_23 sn20_23 78000.000000
Rwneg20_24 in20_24 sn20_24 202000.000000
Rwneg20_25 in20_25 sn20_25 78000.000000
Rwneg20_26 in20_26 sn20_26 78000.000000
Rwneg20_27 in20_27 sn20_27 202000.000000
Rwneg20_28 in20_28 sn20_28 202000.000000
Rwneg20_29 in20_29 sn20_29 78000.000000
Rwneg20_30 in20_30 sn20_30 78000.000000
Rwneg20_31 in20_31 sn20_31 78000.000000
Rwneg20_32 in20_32 sn20_32 202000.000000
Rwneg20_33 in20_33 sn20_33 78000.000000
Rwneg20_34 in20_34 sn20_34 78000.000000
Rwneg20_35 in20_35 sn20_35 202000.000000
Rwneg20_36 in20_36 sn20_36 202000.000000
Rwneg20_37 in20_37 sn20_37 78000.000000
Rwneg20_38 in20_38 sn20_38 202000.000000
Rwneg20_39 in20_39 sn20_39 202000.000000
Rwneg20_40 in20_40 sn20_40 78000.000000
Rwneg20_41 in20_41 sn20_41 78000.000000
Rwneg20_42 in20_42 sn20_42 78000.000000
Rwneg20_43 in20_43 sn20_43 78000.000000
Rwneg20_44 in20_44 sn20_44 78000.000000
Rwneg20_45 in20_45 sn20_45 202000.000000
Rwneg20_46 in20_46 sn20_46 78000.000000
Rwneg20_47 in20_47 sn20_47 78000.000000
Rwneg20_48 in20_48 sn20_48 202000.000000
Rwneg20_49 in20_49 sn20_49 78000.000000
Rwneg20_50 in20_50 sn20_50 78000.000000
Rwneg20_51 in20_51 sn20_51 202000.000000
Rwneg20_52 in20_52 sn20_52 78000.000000
Rwneg20_53 in20_53 sn20_53 78000.000000
Rwneg20_54 in20_54 sn20_54 78000.000000
Rwneg20_55 in20_55 sn20_55 78000.000000
Rwneg20_56 in20_56 sn20_56 202000.000000
Rwneg20_57 in20_57 sn20_57 202000.000000
Rwneg20_58 in20_58 sn20_58 78000.000000
Rwneg20_59 in20_59 sn20_59 202000.000000
Rwneg20_60 in20_60 sn20_60 202000.000000
Rwneg20_61 in20_61 sn20_61 202000.000000
Rwneg20_62 in20_62 sn20_62 78000.000000
Rwneg20_63 in20_63 sn20_63 202000.000000
Rwneg20_64 in20_64 sn20_64 78000.000000
Rwneg20_65 in20_65 sn20_65 202000.000000
Rwneg20_66 in20_66 sn20_66 202000.000000
Rwneg20_67 in20_67 sn20_67 202000.000000
Rwneg20_68 in20_68 sn20_68 202000.000000
Rwneg20_69 in20_69 sn20_69 202000.000000
Rwneg20_70 in20_70 sn20_70 202000.000000
Rwneg20_71 in20_71 sn20_71 202000.000000
Rwneg20_72 in20_72 sn20_72 202000.000000
Rwneg20_73 in20_73 sn20_73 202000.000000
Rwneg20_74 in20_74 sn20_74 202000.000000
Rwneg20_75 in20_75 sn20_75 202000.000000
Rwneg20_76 in20_76 sn20_76 78000.000000
Rwneg20_77 in20_77 sn20_77 78000.000000
Rwneg20_78 in20_78 sn20_78 202000.000000
Rwneg20_79 in20_79 sn20_79 202000.000000
Rwneg20_80 in20_80 sn20_80 78000.000000
Rwneg20_81 in20_81 sn20_81 202000.000000
Rwneg20_82 in20_82 sn20_82 202000.000000
Rwneg20_83 in20_83 sn20_83 202000.000000
Rwneg20_84 in20_84 sn20_84 202000.000000
Rwneg21_1 in21_1 sn21_1 78000.000000
Rwneg21_2 in21_2 sn21_2 202000.000000
Rwneg21_3 in21_3 sn21_3 202000.000000
Rwneg21_4 in21_4 sn21_4 202000.000000
Rwneg21_5 in21_5 sn21_5 202000.000000
Rwneg21_6 in21_6 sn21_6 202000.000000
Rwneg21_7 in21_7 sn21_7 202000.000000
Rwneg21_8 in21_8 sn21_8 202000.000000
Rwneg21_9 in21_9 sn21_9 202000.000000
Rwneg21_10 in21_10 sn21_10 202000.000000
Rwneg21_11 in21_11 sn21_11 78000.000000
Rwneg21_12 in21_12 sn21_12 202000.000000
Rwneg21_13 in21_13 sn21_13 202000.000000
Rwneg21_14 in21_14 sn21_14 202000.000000
Rwneg21_15 in21_15 sn21_15 78000.000000
Rwneg21_16 in21_16 sn21_16 78000.000000
Rwneg21_17 in21_17 sn21_17 78000.000000
Rwneg21_18 in21_18 sn21_18 202000.000000
Rwneg21_19 in21_19 sn21_19 78000.000000
Rwneg21_20 in21_20 sn21_20 78000.000000
Rwneg21_21 in21_21 sn21_21 78000.000000
Rwneg21_22 in21_22 sn21_22 78000.000000
Rwneg21_23 in21_23 sn21_23 78000.000000
Rwneg21_24 in21_24 sn21_24 78000.000000
Rwneg21_25 in21_25 sn21_25 78000.000000
Rwneg21_26 in21_26 sn21_26 78000.000000
Rwneg21_27 in21_27 sn21_27 202000.000000
Rwneg21_28 in21_28 sn21_28 78000.000000
Rwneg21_29 in21_29 sn21_29 78000.000000
Rwneg21_30 in21_30 sn21_30 202000.000000
Rwneg21_31 in21_31 sn21_31 78000.000000
Rwneg21_32 in21_32 sn21_32 202000.000000
Rwneg21_33 in21_33 sn21_33 202000.000000
Rwneg21_34 in21_34 sn21_34 78000.000000
Rwneg21_35 in21_35 sn21_35 202000.000000
Rwneg21_36 in21_36 sn21_36 202000.000000
Rwneg21_37 in21_37 sn21_37 78000.000000
Rwneg21_38 in21_38 sn21_38 78000.000000
Rwneg21_39 in21_39 sn21_39 202000.000000
Rwneg21_40 in21_40 sn21_40 78000.000000
Rwneg21_41 in21_41 sn21_41 202000.000000
Rwneg21_42 in21_42 sn21_42 202000.000000
Rwneg21_43 in21_43 sn21_43 202000.000000
Rwneg21_44 in21_44 sn21_44 202000.000000
Rwneg21_45 in21_45 sn21_45 202000.000000
Rwneg21_46 in21_46 sn21_46 78000.000000
Rwneg21_47 in21_47 sn21_47 202000.000000
Rwneg21_48 in21_48 sn21_48 78000.000000
Rwneg21_49 in21_49 sn21_49 202000.000000
Rwneg21_50 in21_50 sn21_50 202000.000000
Rwneg21_51 in21_51 sn21_51 202000.000000
Rwneg21_52 in21_52 sn21_52 202000.000000
Rwneg21_53 in21_53 sn21_53 78000.000000
Rwneg21_54 in21_54 sn21_54 202000.000000
Rwneg21_55 in21_55 sn21_55 202000.000000
Rwneg21_56 in21_56 sn21_56 202000.000000
Rwneg21_57 in21_57 sn21_57 78000.000000
Rwneg21_58 in21_58 sn21_58 78000.000000
Rwneg21_59 in21_59 sn21_59 202000.000000
Rwneg21_60 in21_60 sn21_60 202000.000000
Rwneg21_61 in21_61 sn21_61 202000.000000
Rwneg21_62 in21_62 sn21_62 78000.000000
Rwneg21_63 in21_63 sn21_63 202000.000000
Rwneg21_64 in21_64 sn21_64 202000.000000
Rwneg21_65 in21_65 sn21_65 202000.000000
Rwneg21_66 in21_66 sn21_66 202000.000000
Rwneg21_67 in21_67 sn21_67 78000.000000
Rwneg21_68 in21_68 sn21_68 202000.000000
Rwneg21_69 in21_69 sn21_69 202000.000000
Rwneg21_70 in21_70 sn21_70 78000.000000
Rwneg21_71 in21_71 sn21_71 202000.000000
Rwneg21_72 in21_72 sn21_72 78000.000000
Rwneg21_73 in21_73 sn21_73 78000.000000
Rwneg21_74 in21_74 sn21_74 78000.000000
Rwneg21_75 in21_75 sn21_75 78000.000000
Rwneg21_76 in21_76 sn21_76 202000.000000
Rwneg21_77 in21_77 sn21_77 78000.000000
Rwneg21_78 in21_78 sn21_78 78000.000000
Rwneg21_79 in21_79 sn21_79 202000.000000
Rwneg21_80 in21_80 sn21_80 202000.000000
Rwneg21_81 in21_81 sn21_81 202000.000000
Rwneg21_82 in21_82 sn21_82 202000.000000
Rwneg21_83 in21_83 sn21_83 202000.000000
Rwneg21_84 in21_84 sn21_84 202000.000000
Rwneg22_1 in22_1 sn22_1 78000.000000
Rwneg22_2 in22_2 sn22_2 78000.000000
Rwneg22_3 in22_3 sn22_3 202000.000000
Rwneg22_4 in22_4 sn22_4 202000.000000
Rwneg22_5 in22_5 sn22_5 202000.000000
Rwneg22_6 in22_6 sn22_6 78000.000000
Rwneg22_7 in22_7 sn22_7 202000.000000
Rwneg22_8 in22_8 sn22_8 202000.000000
Rwneg22_9 in22_9 sn22_9 202000.000000
Rwneg22_10 in22_10 sn22_10 78000.000000
Rwneg22_11 in22_11 sn22_11 78000.000000
Rwneg22_12 in22_12 sn22_12 202000.000000
Rwneg22_13 in22_13 sn22_13 202000.000000
Rwneg22_14 in22_14 sn22_14 202000.000000
Rwneg22_15 in22_15 sn22_15 202000.000000
Rwneg22_16 in22_16 sn22_16 202000.000000
Rwneg22_17 in22_17 sn22_17 78000.000000
Rwneg22_18 in22_18 sn22_18 202000.000000
Rwneg22_19 in22_19 sn22_19 78000.000000
Rwneg22_20 in22_20 sn22_20 202000.000000
Rwneg22_21 in22_21 sn22_21 78000.000000
Rwneg22_22 in22_22 sn22_22 202000.000000
Rwneg22_23 in22_23 sn22_23 202000.000000
Rwneg22_24 in22_24 sn22_24 202000.000000
Rwneg22_25 in22_25 sn22_25 78000.000000
Rwneg22_26 in22_26 sn22_26 202000.000000
Rwneg22_27 in22_27 sn22_27 202000.000000
Rwneg22_28 in22_28 sn22_28 202000.000000
Rwneg22_29 in22_29 sn22_29 78000.000000
Rwneg22_30 in22_30 sn22_30 78000.000000
Rwneg22_31 in22_31 sn22_31 78000.000000
Rwneg22_32 in22_32 sn22_32 202000.000000
Rwneg22_33 in22_33 sn22_33 202000.000000
Rwneg22_34 in22_34 sn22_34 202000.000000
Rwneg22_35 in22_35 sn22_35 202000.000000
Rwneg22_36 in22_36 sn22_36 202000.000000
Rwneg22_37 in22_37 sn22_37 78000.000000
Rwneg22_38 in22_38 sn22_38 202000.000000
Rwneg22_39 in22_39 sn22_39 202000.000000
Rwneg22_40 in22_40 sn22_40 78000.000000
Rwneg22_41 in22_41 sn22_41 78000.000000
Rwneg22_42 in22_42 sn22_42 78000.000000
Rwneg22_43 in22_43 sn22_43 78000.000000
Rwneg22_44 in22_44 sn22_44 78000.000000
Rwneg22_45 in22_45 sn22_45 202000.000000
Rwneg22_46 in22_46 sn22_46 202000.000000
Rwneg22_47 in22_47 sn22_47 202000.000000
Rwneg22_48 in22_48 sn22_48 78000.000000
Rwneg22_49 in22_49 sn22_49 202000.000000
Rwneg22_50 in22_50 sn22_50 202000.000000
Rwneg22_51 in22_51 sn22_51 202000.000000
Rwneg22_52 in22_52 sn22_52 202000.000000
Rwneg22_53 in22_53 sn22_53 78000.000000
Rwneg22_54 in22_54 sn22_54 78000.000000
Rwneg22_55 in22_55 sn22_55 78000.000000
Rwneg22_56 in22_56 sn22_56 78000.000000
Rwneg22_57 in22_57 sn22_57 202000.000000
Rwneg22_58 in22_58 sn22_58 78000.000000
Rwneg22_59 in22_59 sn22_59 202000.000000
Rwneg22_60 in22_60 sn22_60 202000.000000
Rwneg22_61 in22_61 sn22_61 78000.000000
Rwneg22_62 in22_62 sn22_62 78000.000000
Rwneg22_63 in22_63 sn22_63 202000.000000
Rwneg22_64 in22_64 sn22_64 78000.000000
Rwneg22_65 in22_65 sn22_65 78000.000000
Rwneg22_66 in22_66 sn22_66 202000.000000
Rwneg22_67 in22_67 sn22_67 202000.000000
Rwneg22_68 in22_68 sn22_68 78000.000000
Rwneg22_69 in22_69 sn22_69 202000.000000
Rwneg22_70 in22_70 sn22_70 202000.000000
Rwneg22_71 in22_71 sn22_71 78000.000000
Rwneg22_72 in22_72 sn22_72 202000.000000
Rwneg22_73 in22_73 sn22_73 78000.000000
Rwneg22_74 in22_74 sn22_74 202000.000000
Rwneg22_75 in22_75 sn22_75 202000.000000
Rwneg22_76 in22_76 sn22_76 202000.000000
Rwneg22_77 in22_77 sn22_77 78000.000000
Rwneg22_78 in22_78 sn22_78 202000.000000
Rwneg22_79 in22_79 sn22_79 202000.000000
Rwneg22_80 in22_80 sn22_80 78000.000000
Rwneg22_81 in22_81 sn22_81 78000.000000
Rwneg22_82 in22_82 sn22_82 202000.000000
Rwneg22_83 in22_83 sn22_83 78000.000000
Rwneg22_84 in22_84 sn22_84 202000.000000
Rwneg23_1 in23_1 sn23_1 202000.000000
Rwneg23_2 in23_2 sn23_2 78000.000000
Rwneg23_3 in23_3 sn23_3 202000.000000
Rwneg23_4 in23_4 sn23_4 202000.000000
Rwneg23_5 in23_5 sn23_5 78000.000000
Rwneg23_6 in23_6 sn23_6 78000.000000
Rwneg23_7 in23_7 sn23_7 202000.000000
Rwneg23_8 in23_8 sn23_8 78000.000000
Rwneg23_9 in23_9 sn23_9 202000.000000
Rwneg23_10 in23_10 sn23_10 78000.000000
Rwneg23_11 in23_11 sn23_11 78000.000000
Rwneg23_12 in23_12 sn23_12 78000.000000
Rwneg23_13 in23_13 sn23_13 78000.000000
Rwneg23_14 in23_14 sn23_14 78000.000000
Rwneg23_15 in23_15 sn23_15 202000.000000
Rwneg23_16 in23_16 sn23_16 78000.000000
Rwneg23_17 in23_17 sn23_17 202000.000000
Rwneg23_18 in23_18 sn23_18 78000.000000
Rwneg23_19 in23_19 sn23_19 78000.000000
Rwneg23_20 in23_20 sn23_20 78000.000000
Rwneg23_21 in23_21 sn23_21 78000.000000
Rwneg23_22 in23_22 sn23_22 78000.000000
Rwneg23_23 in23_23 sn23_23 202000.000000
Rwneg23_24 in23_24 sn23_24 202000.000000
Rwneg23_25 in23_25 sn23_25 202000.000000
Rwneg23_26 in23_26 sn23_26 78000.000000
Rwneg23_27 in23_27 sn23_27 78000.000000
Rwneg23_28 in23_28 sn23_28 78000.000000
Rwneg23_29 in23_29 sn23_29 78000.000000
Rwneg23_30 in23_30 sn23_30 202000.000000
Rwneg23_31 in23_31 sn23_31 78000.000000
Rwneg23_32 in23_32 sn23_32 78000.000000
Rwneg23_33 in23_33 sn23_33 202000.000000
Rwneg23_34 in23_34 sn23_34 202000.000000
Rwneg23_35 in23_35 sn23_35 78000.000000
Rwneg23_36 in23_36 sn23_36 202000.000000
Rwneg23_37 in23_37 sn23_37 202000.000000
Rwneg23_38 in23_38 sn23_38 78000.000000
Rwneg23_39 in23_39 sn23_39 202000.000000
Rwneg23_40 in23_40 sn23_40 78000.000000
Rwneg23_41 in23_41 sn23_41 78000.000000
Rwneg23_42 in23_42 sn23_42 202000.000000
Rwneg23_43 in23_43 sn23_43 78000.000000
Rwneg23_44 in23_44 sn23_44 202000.000000
Rwneg23_45 in23_45 sn23_45 78000.000000
Rwneg23_46 in23_46 sn23_46 78000.000000
Rwneg23_47 in23_47 sn23_47 202000.000000
Rwneg23_48 in23_48 sn23_48 78000.000000
Rwneg23_49 in23_49 sn23_49 202000.000000
Rwneg23_50 in23_50 sn23_50 202000.000000
Rwneg23_51 in23_51 sn23_51 78000.000000
Rwneg23_52 in23_52 sn23_52 202000.000000
Rwneg23_53 in23_53 sn23_53 78000.000000
Rwneg23_54 in23_54 sn23_54 202000.000000
Rwneg23_55 in23_55 sn23_55 78000.000000
Rwneg23_56 in23_56 sn23_56 78000.000000
Rwneg23_57 in23_57 sn23_57 202000.000000
Rwneg23_58 in23_58 sn23_58 78000.000000
Rwneg23_59 in23_59 sn23_59 202000.000000
Rwneg23_60 in23_60 sn23_60 202000.000000
Rwneg23_61 in23_61 sn23_61 78000.000000
Rwneg23_62 in23_62 sn23_62 202000.000000
Rwneg23_63 in23_63 sn23_63 202000.000000
Rwneg23_64 in23_64 sn23_64 78000.000000
Rwneg23_65 in23_65 sn23_65 78000.000000
Rwneg23_66 in23_66 sn23_66 202000.000000
Rwneg23_67 in23_67 sn23_67 78000.000000
Rwneg23_68 in23_68 sn23_68 202000.000000
Rwneg23_69 in23_69 sn23_69 202000.000000
Rwneg23_70 in23_70 sn23_70 202000.000000
Rwneg23_71 in23_71 sn23_71 202000.000000
Rwneg23_72 in23_72 sn23_72 202000.000000
Rwneg23_73 in23_73 sn23_73 202000.000000
Rwneg23_74 in23_74 sn23_74 202000.000000
Rwneg23_75 in23_75 sn23_75 202000.000000
Rwneg23_76 in23_76 sn23_76 202000.000000
Rwneg23_77 in23_77 sn23_77 78000.000000
Rwneg23_78 in23_78 sn23_78 78000.000000
Rwneg23_79 in23_79 sn23_79 202000.000000
Rwneg23_80 in23_80 sn23_80 78000.000000
Rwneg23_81 in23_81 sn23_81 202000.000000
Rwneg23_82 in23_82 sn23_82 202000.000000
Rwneg23_83 in23_83 sn23_83 78000.000000
Rwneg23_84 in23_84 sn23_84 78000.000000
Rwneg24_1 in24_1 sn24_1 78000.000000
Rwneg24_2 in24_2 sn24_2 202000.000000
Rwneg24_3 in24_3 sn24_3 202000.000000
Rwneg24_4 in24_4 sn24_4 78000.000000
Rwneg24_5 in24_5 sn24_5 78000.000000
Rwneg24_6 in24_6 sn24_6 78000.000000
Rwneg24_7 in24_7 sn24_7 202000.000000
Rwneg24_8 in24_8 sn24_8 78000.000000
Rwneg24_9 in24_9 sn24_9 78000.000000
Rwneg24_10 in24_10 sn24_10 202000.000000
Rwneg24_11 in24_11 sn24_11 78000.000000
Rwneg24_12 in24_12 sn24_12 78000.000000
Rwneg24_13 in24_13 sn24_13 202000.000000
Rwneg24_14 in24_14 sn24_14 78000.000000
Rwneg24_15 in24_15 sn24_15 202000.000000
Rwneg24_16 in24_16 sn24_16 78000.000000
Rwneg24_17 in24_17 sn24_17 78000.000000
Rwneg24_18 in24_18 sn24_18 78000.000000
Rwneg24_19 in24_19 sn24_19 78000.000000
Rwneg24_20 in24_20 sn24_20 202000.000000
Rwneg24_21 in24_21 sn24_21 78000.000000
Rwneg24_22 in24_22 sn24_22 78000.000000
Rwneg24_23 in24_23 sn24_23 78000.000000
Rwneg24_24 in24_24 sn24_24 202000.000000
Rwneg24_25 in24_25 sn24_25 78000.000000
Rwneg24_26 in24_26 sn24_26 202000.000000
Rwneg24_27 in24_27 sn24_27 78000.000000
Rwneg24_28 in24_28 sn24_28 78000.000000
Rwneg24_29 in24_29 sn24_29 78000.000000
Rwneg24_30 in24_30 sn24_30 202000.000000
Rwneg24_31 in24_31 sn24_31 78000.000000
Rwneg24_32 in24_32 sn24_32 78000.000000
Rwneg24_33 in24_33 sn24_33 202000.000000
Rwneg24_34 in24_34 sn24_34 78000.000000
Rwneg24_35 in24_35 sn24_35 202000.000000
Rwneg24_36 in24_36 sn24_36 202000.000000
Rwneg24_37 in24_37 sn24_37 202000.000000
Rwneg24_38 in24_38 sn24_38 78000.000000
Rwneg24_39 in24_39 sn24_39 78000.000000
Rwneg24_40 in24_40 sn24_40 78000.000000
Rwneg24_41 in24_41 sn24_41 78000.000000
Rwneg24_42 in24_42 sn24_42 202000.000000
Rwneg24_43 in24_43 sn24_43 202000.000000
Rwneg24_44 in24_44 sn24_44 202000.000000
Rwneg24_45 in24_45 sn24_45 202000.000000
Rwneg24_46 in24_46 sn24_46 78000.000000
Rwneg24_47 in24_47 sn24_47 202000.000000
Rwneg24_48 in24_48 sn24_48 78000.000000
Rwneg24_49 in24_49 sn24_49 78000.000000
Rwneg24_50 in24_50 sn24_50 202000.000000
Rwneg24_51 in24_51 sn24_51 78000.000000
Rwneg24_52 in24_52 sn24_52 202000.000000
Rwneg24_53 in24_53 sn24_53 78000.000000
Rwneg24_54 in24_54 sn24_54 78000.000000
Rwneg24_55 in24_55 sn24_55 202000.000000
Rwneg24_56 in24_56 sn24_56 78000.000000
Rwneg24_57 in24_57 sn24_57 202000.000000
Rwneg24_58 in24_58 sn24_58 78000.000000
Rwneg24_59 in24_59 sn24_59 78000.000000
Rwneg24_60 in24_60 sn24_60 202000.000000
Rwneg24_61 in24_61 sn24_61 78000.000000
Rwneg24_62 in24_62 sn24_62 78000.000000
Rwneg24_63 in24_63 sn24_63 202000.000000
Rwneg24_64 in24_64 sn24_64 78000.000000
Rwneg24_65 in24_65 sn24_65 78000.000000
Rwneg24_66 in24_66 sn24_66 202000.000000
Rwneg24_67 in24_67 sn24_67 78000.000000
Rwneg24_68 in24_68 sn24_68 78000.000000
Rwneg24_69 in24_69 sn24_69 78000.000000
Rwneg24_70 in24_70 sn24_70 202000.000000
Rwneg24_71 in24_71 sn24_71 78000.000000
Rwneg24_72 in24_72 sn24_72 202000.000000
Rwneg24_73 in24_73 sn24_73 78000.000000
Rwneg24_74 in24_74 sn24_74 78000.000000
Rwneg24_75 in24_75 sn24_75 202000.000000
Rwneg24_76 in24_76 sn24_76 202000.000000
Rwneg24_77 in24_77 sn24_77 78000.000000
Rwneg24_78 in24_78 sn24_78 78000.000000
Rwneg24_79 in24_79 sn24_79 78000.000000
Rwneg24_80 in24_80 sn24_80 78000.000000
Rwneg24_81 in24_81 sn24_81 202000.000000
Rwneg24_82 in24_82 sn24_82 202000.000000
Rwneg24_83 in24_83 sn24_83 202000.000000
Rwneg24_84 in24_84 sn24_84 202000.000000
Rwneg25_1 in25_1 sn25_1 202000.000000
Rwneg25_2 in25_2 sn25_2 78000.000000
Rwneg25_3 in25_3 sn25_3 78000.000000
Rwneg25_4 in25_4 sn25_4 78000.000000
Rwneg25_5 in25_5 sn25_5 202000.000000
Rwneg25_6 in25_6 sn25_6 78000.000000
Rwneg25_7 in25_7 sn25_7 202000.000000
Rwneg25_8 in25_8 sn25_8 78000.000000
Rwneg25_9 in25_9 sn25_9 78000.000000
Rwneg25_10 in25_10 sn25_10 202000.000000
Rwneg25_11 in25_11 sn25_11 202000.000000
Rwneg25_12 in25_12 sn25_12 78000.000000
Rwneg25_13 in25_13 sn25_13 202000.000000
Rwneg25_14 in25_14 sn25_14 78000.000000
Rwneg25_15 in25_15 sn25_15 78000.000000
Rwneg25_16 in25_16 sn25_16 202000.000000
Rwneg25_17 in25_17 sn25_17 202000.000000
Rwneg25_18 in25_18 sn25_18 78000.000000
Rwneg25_19 in25_19 sn25_19 202000.000000
Rwneg25_20 in25_20 sn25_20 202000.000000
Rwneg25_21 in25_21 sn25_21 78000.000000
Rwneg25_22 in25_22 sn25_22 202000.000000
Rwneg25_23 in25_23 sn25_23 78000.000000
Rwneg25_24 in25_24 sn25_24 202000.000000
Rwneg25_25 in25_25 sn25_25 202000.000000
Rwneg25_26 in25_26 sn25_26 202000.000000
Rwneg25_27 in25_27 sn25_27 78000.000000
Rwneg25_28 in25_28 sn25_28 202000.000000
Rwneg25_29 in25_29 sn25_29 202000.000000
Rwneg25_30 in25_30 sn25_30 202000.000000
Rwneg25_31 in25_31 sn25_31 78000.000000
Rwneg25_32 in25_32 sn25_32 202000.000000
Rwneg25_33 in25_33 sn25_33 202000.000000
Rwneg25_34 in25_34 sn25_34 202000.000000
Rwneg25_35 in25_35 sn25_35 78000.000000
Rwneg25_36 in25_36 sn25_36 202000.000000
Rwneg25_37 in25_37 sn25_37 202000.000000
Rwneg25_38 in25_38 sn25_38 202000.000000
Rwneg25_39 in25_39 sn25_39 202000.000000
Rwneg25_40 in25_40 sn25_40 202000.000000
Rwneg25_41 in25_41 sn25_41 202000.000000
Rwneg25_42 in25_42 sn25_42 202000.000000
Rwneg25_43 in25_43 sn25_43 202000.000000
Rwneg25_44 in25_44 sn25_44 202000.000000
Rwneg25_45 in25_45 sn25_45 78000.000000
Rwneg25_46 in25_46 sn25_46 78000.000000
Rwneg25_47 in25_47 sn25_47 202000.000000
Rwneg25_48 in25_48 sn25_48 78000.000000
Rwneg25_49 in25_49 sn25_49 202000.000000
Rwneg25_50 in25_50 sn25_50 202000.000000
Rwneg25_51 in25_51 sn25_51 202000.000000
Rwneg25_52 in25_52 sn25_52 202000.000000
Rwneg25_53 in25_53 sn25_53 78000.000000
Rwneg25_54 in25_54 sn25_54 78000.000000
Rwneg25_55 in25_55 sn25_55 202000.000000
Rwneg25_56 in25_56 sn25_56 78000.000000
Rwneg25_57 in25_57 sn25_57 78000.000000
Rwneg25_58 in25_58 sn25_58 202000.000000
Rwneg25_59 in25_59 sn25_59 202000.000000
Rwneg25_60 in25_60 sn25_60 78000.000000
Rwneg25_61 in25_61 sn25_61 78000.000000
Rwneg25_62 in25_62 sn25_62 202000.000000
Rwneg25_63 in25_63 sn25_63 202000.000000
Rwneg25_64 in25_64 sn25_64 78000.000000
Rwneg25_65 in25_65 sn25_65 202000.000000
Rwneg25_66 in25_66 sn25_66 78000.000000
Rwneg25_67 in25_67 sn25_67 202000.000000
Rwneg25_68 in25_68 sn25_68 78000.000000
Rwneg25_69 in25_69 sn25_69 202000.000000
Rwneg25_70 in25_70 sn25_70 202000.000000
Rwneg25_71 in25_71 sn25_71 202000.000000
Rwneg25_72 in25_72 sn25_72 78000.000000
Rwneg25_73 in25_73 sn25_73 78000.000000
Rwneg25_74 in25_74 sn25_74 78000.000000
Rwneg25_75 in25_75 sn25_75 78000.000000
Rwneg25_76 in25_76 sn25_76 78000.000000
Rwneg25_77 in25_77 sn25_77 202000.000000
Rwneg25_78 in25_78 sn25_78 202000.000000
Rwneg25_79 in25_79 sn25_79 202000.000000
Rwneg25_80 in25_80 sn25_80 78000.000000
Rwneg25_81 in25_81 sn25_81 78000.000000
Rwneg25_82 in25_82 sn25_82 78000.000000
Rwneg25_83 in25_83 sn25_83 78000.000000
Rwneg25_84 in25_84 sn25_84 78000.000000
Rwneg26_1 in26_1 sn26_1 202000.000000
Rwneg26_2 in26_2 sn26_2 78000.000000
Rwneg26_3 in26_3 sn26_3 202000.000000
Rwneg26_4 in26_4 sn26_4 202000.000000
Rwneg26_5 in26_5 sn26_5 202000.000000
Rwneg26_6 in26_6 sn26_6 78000.000000
Rwneg26_7 in26_7 sn26_7 78000.000000
Rwneg26_8 in26_8 sn26_8 78000.000000
Rwneg26_9 in26_9 sn26_9 78000.000000
Rwneg26_10 in26_10 sn26_10 78000.000000
Rwneg26_11 in26_11 sn26_11 78000.000000
Rwneg26_12 in26_12 sn26_12 78000.000000
Rwneg26_13 in26_13 sn26_13 78000.000000
Rwneg26_14 in26_14 sn26_14 202000.000000
Rwneg26_15 in26_15 sn26_15 78000.000000
Rwneg26_16 in26_16 sn26_16 78000.000000
Rwneg26_17 in26_17 sn26_17 202000.000000
Rwneg26_18 in26_18 sn26_18 202000.000000
Rwneg26_19 in26_19 sn26_19 78000.000000
Rwneg26_20 in26_20 sn26_20 78000.000000
Rwneg26_21 in26_21 sn26_21 202000.000000
Rwneg26_22 in26_22 sn26_22 202000.000000
Rwneg26_23 in26_23 sn26_23 78000.000000
Rwneg26_24 in26_24 sn26_24 202000.000000
Rwneg26_25 in26_25 sn26_25 202000.000000
Rwneg26_26 in26_26 sn26_26 202000.000000
Rwneg26_27 in26_27 sn26_27 202000.000000
Rwneg26_28 in26_28 sn26_28 202000.000000
Rwneg26_29 in26_29 sn26_29 202000.000000
Rwneg26_30 in26_30 sn26_30 202000.000000
Rwneg26_31 in26_31 sn26_31 78000.000000
Rwneg26_32 in26_32 sn26_32 78000.000000
Rwneg26_33 in26_33 sn26_33 202000.000000
Rwneg26_34 in26_34 sn26_34 78000.000000
Rwneg26_35 in26_35 sn26_35 202000.000000
Rwneg26_36 in26_36 sn26_36 78000.000000
Rwneg26_37 in26_37 sn26_37 78000.000000
Rwneg26_38 in26_38 sn26_38 78000.000000
Rwneg26_39 in26_39 sn26_39 202000.000000
Rwneg26_40 in26_40 sn26_40 78000.000000
Rwneg26_41 in26_41 sn26_41 202000.000000
Rwneg26_42 in26_42 sn26_42 202000.000000
Rwneg26_43 in26_43 sn26_43 78000.000000
Rwneg26_44 in26_44 sn26_44 202000.000000
Rwneg26_45 in26_45 sn26_45 78000.000000
Rwneg26_46 in26_46 sn26_46 202000.000000
Rwneg26_47 in26_47 sn26_47 78000.000000
Rwneg26_48 in26_48 sn26_48 78000.000000
Rwneg26_49 in26_49 sn26_49 78000.000000
Rwneg26_50 in26_50 sn26_50 202000.000000
Rwneg26_51 in26_51 sn26_51 202000.000000
Rwneg26_52 in26_52 sn26_52 78000.000000
Rwneg26_53 in26_53 sn26_53 202000.000000
Rwneg26_54 in26_54 sn26_54 78000.000000
Rwneg26_55 in26_55 sn26_55 78000.000000
Rwneg26_56 in26_56 sn26_56 78000.000000
Rwneg26_57 in26_57 sn26_57 202000.000000
Rwneg26_58 in26_58 sn26_58 78000.000000
Rwneg26_59 in26_59 sn26_59 202000.000000
Rwneg26_60 in26_60 sn26_60 202000.000000
Rwneg26_61 in26_61 sn26_61 202000.000000
Rwneg26_62 in26_62 sn26_62 202000.000000
Rwneg26_63 in26_63 sn26_63 202000.000000
Rwneg26_64 in26_64 sn26_64 202000.000000
Rwneg26_65 in26_65 sn26_65 78000.000000
Rwneg26_66 in26_66 sn26_66 78000.000000
Rwneg26_67 in26_67 sn26_67 202000.000000
Rwneg26_68 in26_68 sn26_68 78000.000000
Rwneg26_69 in26_69 sn26_69 78000.000000
Rwneg26_70 in26_70 sn26_70 78000.000000
Rwneg26_71 in26_71 sn26_71 78000.000000
Rwneg26_72 in26_72 sn26_72 202000.000000
Rwneg26_73 in26_73 sn26_73 78000.000000
Rwneg26_74 in26_74 sn26_74 202000.000000
Rwneg26_75 in26_75 sn26_75 202000.000000
Rwneg26_76 in26_76 sn26_76 78000.000000
Rwneg26_77 in26_77 sn26_77 78000.000000
Rwneg26_78 in26_78 sn26_78 202000.000000
Rwneg26_79 in26_79 sn26_79 78000.000000
Rwneg26_80 in26_80 sn26_80 202000.000000
Rwneg26_81 in26_81 sn26_81 202000.000000
Rwneg26_82 in26_82 sn26_82 202000.000000
Rwneg26_83 in26_83 sn26_83 202000.000000
Rwneg26_84 in26_84 sn26_84 202000.000000
Rwneg27_1 in27_1 sn27_1 202000.000000
Rwneg27_2 in27_2 sn27_2 202000.000000
Rwneg27_3 in27_3 sn27_3 78000.000000
Rwneg27_4 in27_4 sn27_4 202000.000000
Rwneg27_5 in27_5 sn27_5 78000.000000
Rwneg27_6 in27_6 sn27_6 78000.000000
Rwneg27_7 in27_7 sn27_7 202000.000000
Rwneg27_8 in27_8 sn27_8 78000.000000
Rwneg27_9 in27_9 sn27_9 78000.000000
Rwneg27_10 in27_10 sn27_10 78000.000000
Rwneg27_11 in27_11 sn27_11 202000.000000
Rwneg27_12 in27_12 sn27_12 78000.000000
Rwneg27_13 in27_13 sn27_13 78000.000000
Rwneg27_14 in27_14 sn27_14 78000.000000
Rwneg27_15 in27_15 sn27_15 78000.000000
Rwneg27_16 in27_16 sn27_16 202000.000000
Rwneg27_17 in27_17 sn27_17 202000.000000
Rwneg27_18 in27_18 sn27_18 78000.000000
Rwneg27_19 in27_19 sn27_19 202000.000000
Rwneg27_20 in27_20 sn27_20 78000.000000
Rwneg27_21 in27_21 sn27_21 202000.000000
Rwneg27_22 in27_22 sn27_22 202000.000000
Rwneg27_23 in27_23 sn27_23 78000.000000
Rwneg27_24 in27_24 sn27_24 202000.000000
Rwneg27_25 in27_25 sn27_25 202000.000000
Rwneg27_26 in27_26 sn27_26 78000.000000
Rwneg27_27 in27_27 sn27_27 78000.000000
Rwneg27_28 in27_28 sn27_28 202000.000000
Rwneg27_29 in27_29 sn27_29 78000.000000
Rwneg27_30 in27_30 sn27_30 202000.000000
Rwneg27_31 in27_31 sn27_31 78000.000000
Rwneg27_32 in27_32 sn27_32 78000.000000
Rwneg27_33 in27_33 sn27_33 202000.000000
Rwneg27_34 in27_34 sn27_34 78000.000000
Rwneg27_35 in27_35 sn27_35 78000.000000
Rwneg27_36 in27_36 sn27_36 78000.000000
Rwneg27_37 in27_37 sn27_37 202000.000000
Rwneg27_38 in27_38 sn27_38 202000.000000
Rwneg27_39 in27_39 sn27_39 78000.000000
Rwneg27_40 in27_40 sn27_40 202000.000000
Rwneg27_41 in27_41 sn27_41 78000.000000
Rwneg27_42 in27_42 sn27_42 202000.000000
Rwneg27_43 in27_43 sn27_43 78000.000000
Rwneg27_44 in27_44 sn27_44 202000.000000
Rwneg27_45 in27_45 sn27_45 78000.000000
Rwneg27_46 in27_46 sn27_46 78000.000000
Rwneg27_47 in27_47 sn27_47 78000.000000
Rwneg27_48 in27_48 sn27_48 202000.000000
Rwneg27_49 in27_49 sn27_49 202000.000000
Rwneg27_50 in27_50 sn27_50 202000.000000
Rwneg27_51 in27_51 sn27_51 202000.000000
Rwneg27_52 in27_52 sn27_52 202000.000000
Rwneg27_53 in27_53 sn27_53 78000.000000
Rwneg27_54 in27_54 sn27_54 202000.000000
Rwneg27_55 in27_55 sn27_55 202000.000000
Rwneg27_56 in27_56 sn27_56 78000.000000
Rwneg27_57 in27_57 sn27_57 202000.000000
Rwneg27_58 in27_58 sn27_58 202000.000000
Rwneg27_59 in27_59 sn27_59 202000.000000
Rwneg27_60 in27_60 sn27_60 202000.000000
Rwneg27_61 in27_61 sn27_61 202000.000000
Rwneg27_62 in27_62 sn27_62 202000.000000
Rwneg27_63 in27_63 sn27_63 78000.000000
Rwneg27_64 in27_64 sn27_64 202000.000000
Rwneg27_65 in27_65 sn27_65 78000.000000
Rwneg27_66 in27_66 sn27_66 78000.000000
Rwneg27_67 in27_67 sn27_67 78000.000000
Rwneg27_68 in27_68 sn27_68 78000.000000
Rwneg27_69 in27_69 sn27_69 78000.000000
Rwneg27_70 in27_70 sn27_70 78000.000000
Rwneg27_71 in27_71 sn27_71 78000.000000
Rwneg27_72 in27_72 sn27_72 202000.000000
Rwneg27_73 in27_73 sn27_73 202000.000000
Rwneg27_74 in27_74 sn27_74 202000.000000
Rwneg27_75 in27_75 sn27_75 78000.000000
Rwneg27_76 in27_76 sn27_76 78000.000000
Rwneg27_77 in27_77 sn27_77 78000.000000
Rwneg27_78 in27_78 sn27_78 202000.000000
Rwneg27_79 in27_79 sn27_79 78000.000000
Rwneg27_80 in27_80 sn27_80 78000.000000
Rwneg27_81 in27_81 sn27_81 78000.000000
Rwneg27_82 in27_82 sn27_82 78000.000000
Rwneg27_83 in27_83 sn27_83 78000.000000
Rwneg27_84 in27_84 sn27_84 78000.000000
Rwneg28_1 in28_1 sn28_1 202000.000000
Rwneg28_2 in28_2 sn28_2 78000.000000
Rwneg28_3 in28_3 sn28_3 202000.000000
Rwneg28_4 in28_4 sn28_4 202000.000000
Rwneg28_5 in28_5 sn28_5 202000.000000
Rwneg28_6 in28_6 sn28_6 78000.000000
Rwneg28_7 in28_7 sn28_7 78000.000000
Rwneg28_8 in28_8 sn28_8 202000.000000
Rwneg28_9 in28_9 sn28_9 202000.000000
Rwneg28_10 in28_10 sn28_10 78000.000000
Rwneg28_11 in28_11 sn28_11 78000.000000
Rwneg28_12 in28_12 sn28_12 202000.000000
Rwneg28_13 in28_13 sn28_13 78000.000000
Rwneg28_14 in28_14 sn28_14 202000.000000
Rwneg28_15 in28_15 sn28_15 78000.000000
Rwneg28_16 in28_16 sn28_16 202000.000000
Rwneg28_17 in28_17 sn28_17 78000.000000
Rwneg28_18 in28_18 sn28_18 202000.000000
Rwneg28_19 in28_19 sn28_19 78000.000000
Rwneg28_20 in28_20 sn28_20 78000.000000
Rwneg28_21 in28_21 sn28_21 202000.000000
Rwneg28_22 in28_22 sn28_22 78000.000000
Rwneg28_23 in28_23 sn28_23 78000.000000
Rwneg28_24 in28_24 sn28_24 78000.000000
Rwneg28_25 in28_25 sn28_25 202000.000000
Rwneg28_26 in28_26 sn28_26 202000.000000
Rwneg28_27 in28_27 sn28_27 202000.000000
Rwneg28_28 in28_28 sn28_28 202000.000000
Rwneg28_29 in28_29 sn28_29 78000.000000
Rwneg28_30 in28_30 sn28_30 202000.000000
Rwneg28_31 in28_31 sn28_31 202000.000000
Rwneg28_32 in28_32 sn28_32 78000.000000
Rwneg28_33 in28_33 sn28_33 78000.000000
Rwneg28_34 in28_34 sn28_34 202000.000000
Rwneg28_35 in28_35 sn28_35 202000.000000
Rwneg28_36 in28_36 sn28_36 202000.000000
Rwneg28_37 in28_37 sn28_37 202000.000000
Rwneg28_38 in28_38 sn28_38 202000.000000
Rwneg28_39 in28_39 sn28_39 202000.000000
Rwneg28_40 in28_40 sn28_40 78000.000000
Rwneg28_41 in28_41 sn28_41 202000.000000
Rwneg28_42 in28_42 sn28_42 202000.000000
Rwneg28_43 in28_43 sn28_43 202000.000000
Rwneg28_44 in28_44 sn28_44 202000.000000
Rwneg28_45 in28_45 sn28_45 78000.000000
Rwneg28_46 in28_46 sn28_46 202000.000000
Rwneg28_47 in28_47 sn28_47 202000.000000
Rwneg28_48 in28_48 sn28_48 78000.000000
Rwneg28_49 in28_49 sn28_49 202000.000000
Rwneg28_50 in28_50 sn28_50 202000.000000
Rwneg28_51 in28_51 sn28_51 202000.000000
Rwneg28_52 in28_52 sn28_52 202000.000000
Rwneg28_53 in28_53 sn28_53 78000.000000
Rwneg28_54 in28_54 sn28_54 202000.000000
Rwneg28_55 in28_55 sn28_55 78000.000000
Rwneg28_56 in28_56 sn28_56 202000.000000
Rwneg28_57 in28_57 sn28_57 202000.000000
Rwneg28_58 in28_58 sn28_58 78000.000000
Rwneg28_59 in28_59 sn28_59 202000.000000
Rwneg28_60 in28_60 sn28_60 202000.000000
Rwneg28_61 in28_61 sn28_61 202000.000000
Rwneg28_62 in28_62 sn28_62 78000.000000
Rwneg28_63 in28_63 sn28_63 202000.000000
Rwneg28_64 in28_64 sn28_64 78000.000000
Rwneg28_65 in28_65 sn28_65 78000.000000
Rwneg28_66 in28_66 sn28_66 202000.000000
Rwneg28_67 in28_67 sn28_67 202000.000000
Rwneg28_68 in28_68 sn28_68 202000.000000
Rwneg28_69 in28_69 sn28_69 202000.000000
Rwneg28_70 in28_70 sn28_70 78000.000000
Rwneg28_71 in28_71 sn28_71 78000.000000
Rwneg28_72 in28_72 sn28_72 202000.000000
Rwneg28_73 in28_73 sn28_73 202000.000000
Rwneg28_74 in28_74 sn28_74 202000.000000
Rwneg28_75 in28_75 sn28_75 202000.000000
Rwneg28_76 in28_76 sn28_76 202000.000000
Rwneg28_77 in28_77 sn28_77 78000.000000
Rwneg28_78 in28_78 sn28_78 202000.000000
Rwneg28_79 in28_79 sn28_79 202000.000000
Rwneg28_80 in28_80 sn28_80 78000.000000
Rwneg28_81 in28_81 sn28_81 78000.000000
Rwneg28_82 in28_82 sn28_82 202000.000000
Rwneg28_83 in28_83 sn28_83 202000.000000
Rwneg28_84 in28_84 sn28_84 78000.000000
Rwneg29_1 in29_1 sn29_1 78000.000000
Rwneg29_2 in29_2 sn29_2 202000.000000
Rwneg29_3 in29_3 sn29_3 78000.000000
Rwneg29_4 in29_4 sn29_4 78000.000000
Rwneg29_5 in29_5 sn29_5 78000.000000
Rwneg29_6 in29_6 sn29_6 202000.000000
Rwneg29_7 in29_7 sn29_7 78000.000000
Rwneg29_8 in29_8 sn29_8 202000.000000
Rwneg29_9 in29_9 sn29_9 78000.000000
Rwneg29_10 in29_10 sn29_10 78000.000000
Rwneg29_11 in29_11 sn29_11 202000.000000
Rwneg29_12 in29_12 sn29_12 202000.000000
Rwneg29_13 in29_13 sn29_13 202000.000000
Rwneg29_14 in29_14 sn29_14 78000.000000
Rwneg29_15 in29_15 sn29_15 202000.000000
Rwneg29_16 in29_16 sn29_16 202000.000000
Rwneg29_17 in29_17 sn29_17 202000.000000
Rwneg29_18 in29_18 sn29_18 202000.000000
Rwneg29_19 in29_19 sn29_19 202000.000000
Rwneg29_20 in29_20 sn29_20 78000.000000
Rwneg29_21 in29_21 sn29_21 202000.000000
Rwneg29_22 in29_22 sn29_22 202000.000000
Rwneg29_23 in29_23 sn29_23 202000.000000
Rwneg29_24 in29_24 sn29_24 202000.000000
Rwneg29_25 in29_25 sn29_25 78000.000000
Rwneg29_26 in29_26 sn29_26 78000.000000
Rwneg29_27 in29_27 sn29_27 78000.000000
Rwneg29_28 in29_28 sn29_28 78000.000000
Rwneg29_29 in29_29 sn29_29 202000.000000
Rwneg29_30 in29_30 sn29_30 202000.000000
Rwneg29_31 in29_31 sn29_31 202000.000000
Rwneg29_32 in29_32 sn29_32 78000.000000
Rwneg29_33 in29_33 sn29_33 202000.000000
Rwneg29_34 in29_34 sn29_34 78000.000000
Rwneg29_35 in29_35 sn29_35 78000.000000
Rwneg29_36 in29_36 sn29_36 78000.000000
Rwneg29_37 in29_37 sn29_37 78000.000000
Rwneg29_38 in29_38 sn29_38 78000.000000
Rwneg29_39 in29_39 sn29_39 202000.000000
Rwneg29_40 in29_40 sn29_40 78000.000000
Rwneg29_41 in29_41 sn29_41 78000.000000
Rwneg29_42 in29_42 sn29_42 202000.000000
Rwneg29_43 in29_43 sn29_43 78000.000000
Rwneg29_44 in29_44 sn29_44 202000.000000
Rwneg29_45 in29_45 sn29_45 202000.000000
Rwneg29_46 in29_46 sn29_46 78000.000000
Rwneg29_47 in29_47 sn29_47 202000.000000
Rwneg29_48 in29_48 sn29_48 202000.000000
Rwneg29_49 in29_49 sn29_49 78000.000000
Rwneg29_50 in29_50 sn29_50 78000.000000
Rwneg29_51 in29_51 sn29_51 202000.000000
Rwneg29_52 in29_52 sn29_52 78000.000000
Rwneg29_53 in29_53 sn29_53 78000.000000
Rwneg29_54 in29_54 sn29_54 202000.000000
Rwneg29_55 in29_55 sn29_55 202000.000000
Rwneg29_56 in29_56 sn29_56 78000.000000
Rwneg29_57 in29_57 sn29_57 202000.000000
Rwneg29_58 in29_58 sn29_58 78000.000000
Rwneg29_59 in29_59 sn29_59 78000.000000
Rwneg29_60 in29_60 sn29_60 202000.000000
Rwneg29_61 in29_61 sn29_61 202000.000000
Rwneg29_62 in29_62 sn29_62 202000.000000
Rwneg29_63 in29_63 sn29_63 78000.000000
Rwneg29_64 in29_64 sn29_64 202000.000000
Rwneg29_65 in29_65 sn29_65 202000.000000
Rwneg29_66 in29_66 sn29_66 202000.000000
Rwneg29_67 in29_67 sn29_67 78000.000000
Rwneg29_68 in29_68 sn29_68 202000.000000
Rwneg29_69 in29_69 sn29_69 78000.000000
Rwneg29_70 in29_70 sn29_70 202000.000000
Rwneg29_71 in29_71 sn29_71 78000.000000
Rwneg29_72 in29_72 sn29_72 78000.000000
Rwneg29_73 in29_73 sn29_73 202000.000000
Rwneg29_74 in29_74 sn29_74 78000.000000
Rwneg29_75 in29_75 sn29_75 78000.000000
Rwneg29_76 in29_76 sn29_76 78000.000000
Rwneg29_77 in29_77 sn29_77 78000.000000
Rwneg29_78 in29_78 sn29_78 202000.000000
Rwneg29_79 in29_79 sn29_79 78000.000000
Rwneg29_80 in29_80 sn29_80 78000.000000
Rwneg29_81 in29_81 sn29_81 202000.000000
Rwneg29_82 in29_82 sn29_82 78000.000000
Rwneg29_83 in29_83 sn29_83 202000.000000
Rwneg29_84 in29_84 sn29_84 202000.000000
Rwneg30_1 in30_1 sn30_1 202000.000000
Rwneg30_2 in30_2 sn30_2 202000.000000
Rwneg30_3 in30_3 sn30_3 78000.000000
Rwneg30_4 in30_4 sn30_4 78000.000000
Rwneg30_5 in30_5 sn30_5 78000.000000
Rwneg30_6 in30_6 sn30_6 202000.000000
Rwneg30_7 in30_7 sn30_7 78000.000000
Rwneg30_8 in30_8 sn30_8 202000.000000
Rwneg30_9 in30_9 sn30_9 78000.000000
Rwneg30_10 in30_10 sn30_10 202000.000000
Rwneg30_11 in30_11 sn30_11 78000.000000
Rwneg30_12 in30_12 sn30_12 202000.000000
Rwneg30_13 in30_13 sn30_13 202000.000000
Rwneg30_14 in30_14 sn30_14 78000.000000
Rwneg30_15 in30_15 sn30_15 202000.000000
Rwneg30_16 in30_16 sn30_16 202000.000000
Rwneg30_17 in30_17 sn30_17 78000.000000
Rwneg30_18 in30_18 sn30_18 202000.000000
Rwneg30_19 in30_19 sn30_19 202000.000000
Rwneg30_20 in30_20 sn30_20 202000.000000
Rwneg30_21 in30_21 sn30_21 202000.000000
Rwneg30_22 in30_22 sn30_22 202000.000000
Rwneg30_23 in30_23 sn30_23 78000.000000
Rwneg30_24 in30_24 sn30_24 202000.000000
Rwneg30_25 in30_25 sn30_25 202000.000000
Rwneg30_26 in30_26 sn30_26 202000.000000
Rwneg30_27 in30_27 sn30_27 78000.000000
Rwneg30_28 in30_28 sn30_28 202000.000000
Rwneg30_29 in30_29 sn30_29 202000.000000
Rwneg30_30 in30_30 sn30_30 202000.000000
Rwneg30_31 in30_31 sn30_31 78000.000000
Rwneg30_32 in30_32 sn30_32 78000.000000
Rwneg30_33 in30_33 sn30_33 202000.000000
Rwneg30_34 in30_34 sn30_34 78000.000000
Rwneg30_35 in30_35 sn30_35 78000.000000
Rwneg30_36 in30_36 sn30_36 202000.000000
Rwneg30_37 in30_37 sn30_37 78000.000000
Rwneg30_38 in30_38 sn30_38 202000.000000
Rwneg30_39 in30_39 sn30_39 202000.000000
Rwneg30_40 in30_40 sn30_40 202000.000000
Rwneg30_41 in30_41 sn30_41 78000.000000
Rwneg30_42 in30_42 sn30_42 78000.000000
Rwneg30_43 in30_43 sn30_43 78000.000000
Rwneg30_44 in30_44 sn30_44 202000.000000
Rwneg30_45 in30_45 sn30_45 202000.000000
Rwneg30_46 in30_46 sn30_46 78000.000000
Rwneg30_47 in30_47 sn30_47 202000.000000
Rwneg30_48 in30_48 sn30_48 78000.000000
Rwneg30_49 in30_49 sn30_49 202000.000000
Rwneg30_50 in30_50 sn30_50 202000.000000
Rwneg30_51 in30_51 sn30_51 202000.000000
Rwneg30_52 in30_52 sn30_52 78000.000000
Rwneg30_53 in30_53 sn30_53 78000.000000
Rwneg30_54 in30_54 sn30_54 78000.000000
Rwneg30_55 in30_55 sn30_55 202000.000000
Rwneg30_56 in30_56 sn30_56 78000.000000
Rwneg30_57 in30_57 sn30_57 78000.000000
Rwneg30_58 in30_58 sn30_58 78000.000000
Rwneg30_59 in30_59 sn30_59 78000.000000
Rwneg30_60 in30_60 sn30_60 202000.000000
Rwneg30_61 in30_61 sn30_61 202000.000000
Rwneg30_62 in30_62 sn30_62 78000.000000
Rwneg30_63 in30_63 sn30_63 202000.000000
Rwneg30_64 in30_64 sn30_64 78000.000000
Rwneg30_65 in30_65 sn30_65 78000.000000
Rwneg30_66 in30_66 sn30_66 202000.000000
Rwneg30_67 in30_67 sn30_67 202000.000000
Rwneg30_68 in30_68 sn30_68 202000.000000
Rwneg30_69 in30_69 sn30_69 78000.000000
Rwneg30_70 in30_70 sn30_70 78000.000000
Rwneg30_71 in30_71 sn30_71 78000.000000
Rwneg30_72 in30_72 sn30_72 202000.000000
Rwneg30_73 in30_73 sn30_73 78000.000000
Rwneg30_74 in30_74 sn30_74 202000.000000
Rwneg30_75 in30_75 sn30_75 202000.000000
Rwneg30_76 in30_76 sn30_76 78000.000000
Rwneg30_77 in30_77 sn30_77 78000.000000
Rwneg30_78 in30_78 sn30_78 78000.000000
Rwneg30_79 in30_79 sn30_79 78000.000000
Rwneg30_80 in30_80 sn30_80 78000.000000
Rwneg30_81 in30_81 sn30_81 202000.000000
Rwneg30_82 in30_82 sn30_82 202000.000000
Rwneg30_83 in30_83 sn30_83 202000.000000
Rwneg30_84 in30_84 sn30_84 78000.000000
Rwneg31_1 in31_1 sn31_1 202000.000000
Rwneg31_2 in31_2 sn31_2 78000.000000
Rwneg31_3 in31_3 sn31_3 202000.000000
Rwneg31_4 in31_4 sn31_4 202000.000000
Rwneg31_5 in31_5 sn31_5 202000.000000
Rwneg31_6 in31_6 sn31_6 78000.000000
Rwneg31_7 in31_7 sn31_7 78000.000000
Rwneg31_8 in31_8 sn31_8 202000.000000
Rwneg31_9 in31_9 sn31_9 202000.000000
Rwneg31_10 in31_10 sn31_10 202000.000000
Rwneg31_11 in31_11 sn31_11 202000.000000
Rwneg31_12 in31_12 sn31_12 202000.000000
Rwneg31_13 in31_13 sn31_13 202000.000000
Rwneg31_14 in31_14 sn31_14 78000.000000
Rwneg31_15 in31_15 sn31_15 202000.000000
Rwneg31_16 in31_16 sn31_16 78000.000000
Rwneg31_17 in31_17 sn31_17 202000.000000
Rwneg31_18 in31_18 sn31_18 202000.000000
Rwneg31_19 in31_19 sn31_19 78000.000000
Rwneg31_20 in31_20 sn31_20 78000.000000
Rwneg31_21 in31_21 sn31_21 78000.000000
Rwneg31_22 in31_22 sn31_22 202000.000000
Rwneg31_23 in31_23 sn31_23 202000.000000
Rwneg31_24 in31_24 sn31_24 202000.000000
Rwneg31_25 in31_25 sn31_25 202000.000000
Rwneg31_26 in31_26 sn31_26 202000.000000
Rwneg31_27 in31_27 sn31_27 202000.000000
Rwneg31_28 in31_28 sn31_28 78000.000000
Rwneg31_29 in31_29 sn31_29 78000.000000
Rwneg31_30 in31_30 sn31_30 78000.000000
Rwneg31_31 in31_31 sn31_31 202000.000000
Rwneg31_32 in31_32 sn31_32 202000.000000
Rwneg31_33 in31_33 sn31_33 78000.000000
Rwneg31_34 in31_34 sn31_34 202000.000000
Rwneg31_35 in31_35 sn31_35 78000.000000
Rwneg31_36 in31_36 sn31_36 202000.000000
Rwneg31_37 in31_37 sn31_37 78000.000000
Rwneg31_38 in31_38 sn31_38 78000.000000
Rwneg31_39 in31_39 sn31_39 202000.000000
Rwneg31_40 in31_40 sn31_40 78000.000000
Rwneg31_41 in31_41 sn31_41 202000.000000
Rwneg31_42 in31_42 sn31_42 78000.000000
Rwneg31_43 in31_43 sn31_43 78000.000000
Rwneg31_44 in31_44 sn31_44 202000.000000
Rwneg31_45 in31_45 sn31_45 78000.000000
Rwneg31_46 in31_46 sn31_46 78000.000000
Rwneg31_47 in31_47 sn31_47 202000.000000
Rwneg31_48 in31_48 sn31_48 78000.000000
Rwneg31_49 in31_49 sn31_49 202000.000000
Rwneg31_50 in31_50 sn31_50 78000.000000
Rwneg31_51 in31_51 sn31_51 78000.000000
Rwneg31_52 in31_52 sn31_52 78000.000000
Rwneg31_53 in31_53 sn31_53 202000.000000
Rwneg31_54 in31_54 sn31_54 202000.000000
Rwneg31_55 in31_55 sn31_55 78000.000000
Rwneg31_56 in31_56 sn31_56 202000.000000
Rwneg31_57 in31_57 sn31_57 202000.000000
Rwneg31_58 in31_58 sn31_58 202000.000000
Rwneg31_59 in31_59 sn31_59 202000.000000
Rwneg31_60 in31_60 sn31_60 202000.000000
Rwneg31_61 in31_61 sn31_61 202000.000000
Rwneg31_62 in31_62 sn31_62 202000.000000
Rwneg31_63 in31_63 sn31_63 202000.000000
Rwneg31_64 in31_64 sn31_64 78000.000000
Rwneg31_65 in31_65 sn31_65 202000.000000
Rwneg31_66 in31_66 sn31_66 202000.000000
Rwneg31_67 in31_67 sn31_67 78000.000000
Rwneg31_68 in31_68 sn31_68 202000.000000
Rwneg31_69 in31_69 sn31_69 202000.000000
Rwneg31_70 in31_70 sn31_70 78000.000000
Rwneg31_71 in31_71 sn31_71 202000.000000
Rwneg31_72 in31_72 sn31_72 202000.000000
Rwneg31_73 in31_73 sn31_73 202000.000000
Rwneg31_74 in31_74 sn31_74 78000.000000
Rwneg31_75 in31_75 sn31_75 78000.000000
Rwneg31_76 in31_76 sn31_76 202000.000000
Rwneg31_77 in31_77 sn31_77 78000.000000
Rwneg31_78 in31_78 sn31_78 202000.000000
Rwneg31_79 in31_79 sn31_79 202000.000000
Rwneg31_80 in31_80 sn31_80 202000.000000
Rwneg31_81 in31_81 sn31_81 202000.000000
Rwneg31_82 in31_82 sn31_82 202000.000000
Rwneg31_83 in31_83 sn31_83 202000.000000
Rwneg31_84 in31_84 sn31_84 78000.000000
Rwneg32_1 in32_1 sn32_1 78000.000000
Rwneg32_2 in32_2 sn32_2 78000.000000
Rwneg32_3 in32_3 sn32_3 78000.000000
Rwneg32_4 in32_4 sn32_4 202000.000000
Rwneg32_5 in32_5 sn32_5 202000.000000
Rwneg32_6 in32_6 sn32_6 202000.000000
Rwneg32_7 in32_7 sn32_7 78000.000000
Rwneg32_8 in32_8 sn32_8 202000.000000
Rwneg32_9 in32_9 sn32_9 202000.000000
Rwneg32_10 in32_10 sn32_10 78000.000000
Rwneg32_11 in32_11 sn32_11 202000.000000
Rwneg32_12 in32_12 sn32_12 78000.000000
Rwneg32_13 in32_13 sn32_13 202000.000000
Rwneg32_14 in32_14 sn32_14 202000.000000
Rwneg32_15 in32_15 sn32_15 202000.000000
Rwneg32_16 in32_16 sn32_16 202000.000000
Rwneg32_17 in32_17 sn32_17 202000.000000
Rwneg32_18 in32_18 sn32_18 78000.000000
Rwneg32_19 in32_19 sn32_19 202000.000000
Rwneg32_20 in32_20 sn32_20 78000.000000
Rwneg32_21 in32_21 sn32_21 202000.000000
Rwneg32_22 in32_22 sn32_22 202000.000000
Rwneg32_23 in32_23 sn32_23 202000.000000
Rwneg32_24 in32_24 sn32_24 78000.000000
Rwneg32_25 in32_25 sn32_25 78000.000000
Rwneg32_26 in32_26 sn32_26 202000.000000
Rwneg32_27 in32_27 sn32_27 202000.000000
Rwneg32_28 in32_28 sn32_28 78000.000000
Rwneg32_29 in32_29 sn32_29 78000.000000
Rwneg32_30 in32_30 sn32_30 202000.000000
Rwneg32_31 in32_31 sn32_31 202000.000000
Rwneg32_32 in32_32 sn32_32 202000.000000
Rwneg32_33 in32_33 sn32_33 78000.000000
Rwneg32_34 in32_34 sn32_34 78000.000000
Rwneg32_35 in32_35 sn32_35 202000.000000
Rwneg32_36 in32_36 sn32_36 78000.000000
Rwneg32_37 in32_37 sn32_37 202000.000000
Rwneg32_38 in32_38 sn32_38 78000.000000
Rwneg32_39 in32_39 sn32_39 202000.000000
Rwneg32_40 in32_40 sn32_40 202000.000000
Rwneg32_41 in32_41 sn32_41 78000.000000
Rwneg32_42 in32_42 sn32_42 202000.000000
Rwneg32_43 in32_43 sn32_43 202000.000000
Rwneg32_44 in32_44 sn32_44 78000.000000
Rwneg32_45 in32_45 sn32_45 78000.000000
Rwneg32_46 in32_46 sn32_46 202000.000000
Rwneg32_47 in32_47 sn32_47 78000.000000
Rwneg32_48 in32_48 sn32_48 78000.000000
Rwneg32_49 in32_49 sn32_49 78000.000000
Rwneg32_50 in32_50 sn32_50 78000.000000
Rwneg32_51 in32_51 sn32_51 78000.000000
Rwneg32_52 in32_52 sn32_52 78000.000000
Rwneg32_53 in32_53 sn32_53 78000.000000
Rwneg32_54 in32_54 sn32_54 202000.000000
Rwneg32_55 in32_55 sn32_55 78000.000000
Rwneg32_56 in32_56 sn32_56 78000.000000
Rwneg32_57 in32_57 sn32_57 78000.000000
Rwneg32_58 in32_58 sn32_58 202000.000000
Rwneg32_59 in32_59 sn32_59 202000.000000
Rwneg32_60 in32_60 sn32_60 78000.000000
Rwneg32_61 in32_61 sn32_61 78000.000000
Rwneg32_62 in32_62 sn32_62 202000.000000
Rwneg32_63 in32_63 sn32_63 202000.000000
Rwneg32_64 in32_64 sn32_64 78000.000000
Rwneg32_65 in32_65 sn32_65 78000.000000
Rwneg32_66 in32_66 sn32_66 78000.000000
Rwneg32_67 in32_67 sn32_67 202000.000000
Rwneg32_68 in32_68 sn32_68 78000.000000
Rwneg32_69 in32_69 sn32_69 202000.000000
Rwneg32_70 in32_70 sn32_70 202000.000000
Rwneg32_71 in32_71 sn32_71 78000.000000
Rwneg32_72 in32_72 sn32_72 78000.000000
Rwneg32_73 in32_73 sn32_73 78000.000000
Rwneg32_74 in32_74 sn32_74 78000.000000
Rwneg32_75 in32_75 sn32_75 78000.000000
Rwneg32_76 in32_76 sn32_76 78000.000000
Rwneg32_77 in32_77 sn32_77 202000.000000
Rwneg32_78 in32_78 sn32_78 202000.000000
Rwneg32_79 in32_79 sn32_79 202000.000000
Rwneg32_80 in32_80 sn32_80 202000.000000
Rwneg32_81 in32_81 sn32_81 202000.000000
Rwneg32_82 in32_82 sn32_82 78000.000000
Rwneg32_83 in32_83 sn32_83 202000.000000
Rwneg32_84 in32_84 sn32_84 202000.000000
Rwneg33_1 in33_1 sn33_1 78000.000000
Rwneg33_2 in33_2 sn33_2 78000.000000
Rwneg33_3 in33_3 sn33_3 202000.000000
Rwneg33_4 in33_4 sn33_4 202000.000000
Rwneg33_5 in33_5 sn33_5 202000.000000
Rwneg33_6 in33_6 sn33_6 202000.000000
Rwneg33_7 in33_7 sn33_7 78000.000000
Rwneg33_8 in33_8 sn33_8 202000.000000
Rwneg33_9 in33_9 sn33_9 78000.000000
Rwneg33_10 in33_10 sn33_10 78000.000000
Rwneg33_11 in33_11 sn33_11 78000.000000
Rwneg33_12 in33_12 sn33_12 202000.000000
Rwneg33_13 in33_13 sn33_13 202000.000000
Rwneg33_14 in33_14 sn33_14 78000.000000
Rwneg33_15 in33_15 sn33_15 202000.000000
Rwneg33_16 in33_16 sn33_16 78000.000000
Rwneg33_17 in33_17 sn33_17 202000.000000
Rwneg33_18 in33_18 sn33_18 202000.000000
Rwneg33_19 in33_19 sn33_19 202000.000000
Rwneg33_20 in33_20 sn33_20 202000.000000
Rwneg33_21 in33_21 sn33_21 202000.000000
Rwneg33_22 in33_22 sn33_22 202000.000000
Rwneg33_23 in33_23 sn33_23 202000.000000
Rwneg33_24 in33_24 sn33_24 202000.000000
Rwneg33_25 in33_25 sn33_25 202000.000000
Rwneg33_26 in33_26 sn33_26 78000.000000
Rwneg33_27 in33_27 sn33_27 78000.000000
Rwneg33_28 in33_28 sn33_28 202000.000000
Rwneg33_29 in33_29 sn33_29 78000.000000
Rwneg33_30 in33_30 sn33_30 202000.000000
Rwneg33_31 in33_31 sn33_31 78000.000000
Rwneg33_32 in33_32 sn33_32 78000.000000
Rwneg33_33 in33_33 sn33_33 202000.000000
Rwneg33_34 in33_34 sn33_34 78000.000000
Rwneg33_35 in33_35 sn33_35 78000.000000
Rwneg33_36 in33_36 sn33_36 202000.000000
Rwneg33_37 in33_37 sn33_37 78000.000000
Rwneg33_38 in33_38 sn33_38 202000.000000
Rwneg33_39 in33_39 sn33_39 202000.000000
Rwneg33_40 in33_40 sn33_40 202000.000000
Rwneg33_41 in33_41 sn33_41 202000.000000
Rwneg33_42 in33_42 sn33_42 78000.000000
Rwneg33_43 in33_43 sn33_43 202000.000000
Rwneg33_44 in33_44 sn33_44 202000.000000
Rwneg33_45 in33_45 sn33_45 202000.000000
Rwneg33_46 in33_46 sn33_46 78000.000000
Rwneg33_47 in33_47 sn33_47 202000.000000
Rwneg33_48 in33_48 sn33_48 202000.000000
Rwneg33_49 in33_49 sn33_49 78000.000000
Rwneg33_50 in33_50 sn33_50 78000.000000
Rwneg33_51 in33_51 sn33_51 78000.000000
Rwneg33_52 in33_52 sn33_52 78000.000000
Rwneg33_53 in33_53 sn33_53 202000.000000
Rwneg33_54 in33_54 sn33_54 202000.000000
Rwneg33_55 in33_55 sn33_55 78000.000000
Rwneg33_56 in33_56 sn33_56 78000.000000
Rwneg33_57 in33_57 sn33_57 202000.000000
Rwneg33_58 in33_58 sn33_58 202000.000000
Rwneg33_59 in33_59 sn33_59 78000.000000
Rwneg33_60 in33_60 sn33_60 202000.000000
Rwneg33_61 in33_61 sn33_61 202000.000000
Rwneg33_62 in33_62 sn33_62 202000.000000
Rwneg33_63 in33_63 sn33_63 202000.000000
Rwneg33_64 in33_64 sn33_64 202000.000000
Rwneg33_65 in33_65 sn33_65 78000.000000
Rwneg33_66 in33_66 sn33_66 202000.000000
Rwneg33_67 in33_67 sn33_67 202000.000000
Rwneg33_68 in33_68 sn33_68 202000.000000
Rwneg33_69 in33_69 sn33_69 78000.000000
Rwneg33_70 in33_70 sn33_70 202000.000000
Rwneg33_71 in33_71 sn33_71 202000.000000
Rwneg33_72 in33_72 sn33_72 78000.000000
Rwneg33_73 in33_73 sn33_73 78000.000000
Rwneg33_74 in33_74 sn33_74 78000.000000
Rwneg33_75 in33_75 sn33_75 202000.000000
Rwneg33_76 in33_76 sn33_76 78000.000000
Rwneg33_77 in33_77 sn33_77 202000.000000
Rwneg33_78 in33_78 sn33_78 78000.000000
Rwneg33_79 in33_79 sn33_79 202000.000000
Rwneg33_80 in33_80 sn33_80 78000.000000
Rwneg33_81 in33_81 sn33_81 202000.000000
Rwneg33_82 in33_82 sn33_82 78000.000000
Rwneg33_83 in33_83 sn33_83 202000.000000
Rwneg33_84 in33_84 sn33_84 202000.000000
Rwneg34_1 in34_1 sn34_1 202000.000000
Rwneg34_2 in34_2 sn34_2 78000.000000
Rwneg34_3 in34_3 sn34_3 78000.000000
Rwneg34_4 in34_4 sn34_4 78000.000000
Rwneg34_5 in34_5 sn34_5 78000.000000
Rwneg34_6 in34_6 sn34_6 202000.000000
Rwneg34_7 in34_7 sn34_7 78000.000000
Rwneg34_8 in34_8 sn34_8 78000.000000
Rwneg34_9 in34_9 sn34_9 78000.000000
Rwneg34_10 in34_10 sn34_10 202000.000000
Rwneg34_11 in34_11 sn34_11 202000.000000
Rwneg34_12 in34_12 sn34_12 202000.000000
Rwneg34_13 in34_13 sn34_13 202000.000000
Rwneg34_14 in34_14 sn34_14 78000.000000
Rwneg34_15 in34_15 sn34_15 202000.000000
Rwneg34_16 in34_16 sn34_16 202000.000000
Rwneg34_17 in34_17 sn34_17 78000.000000
Rwneg34_18 in34_18 sn34_18 202000.000000
Rwneg34_19 in34_19 sn34_19 202000.000000
Rwneg34_20 in34_20 sn34_20 202000.000000
Rwneg34_21 in34_21 sn34_21 202000.000000
Rwneg34_22 in34_22 sn34_22 202000.000000
Rwneg34_23 in34_23 sn34_23 78000.000000
Rwneg34_24 in34_24 sn34_24 202000.000000
Rwneg34_25 in34_25 sn34_25 202000.000000
Rwneg34_26 in34_26 sn34_26 202000.000000
Rwneg34_27 in34_27 sn34_27 78000.000000
Rwneg34_28 in34_28 sn34_28 202000.000000
Rwneg34_29 in34_29 sn34_29 78000.000000
Rwneg34_30 in34_30 sn34_30 202000.000000
Rwneg34_31 in34_31 sn34_31 78000.000000
Rwneg34_32 in34_32 sn34_32 202000.000000
Rwneg34_33 in34_33 sn34_33 202000.000000
Rwneg34_34 in34_34 sn34_34 202000.000000
Rwneg34_35 in34_35 sn34_35 78000.000000
Rwneg34_36 in34_36 sn34_36 202000.000000
Rwneg34_37 in34_37 sn34_37 78000.000000
Rwneg34_38 in34_38 sn34_38 202000.000000
Rwneg34_39 in34_39 sn34_39 202000.000000
Rwneg34_40 in34_40 sn34_40 202000.000000
Rwneg34_41 in34_41 sn34_41 78000.000000
Rwneg34_42 in34_42 sn34_42 78000.000000
Rwneg34_43 in34_43 sn34_43 78000.000000
Rwneg34_44 in34_44 sn34_44 202000.000000
Rwneg34_45 in34_45 sn34_45 202000.000000
Rwneg34_46 in34_46 sn34_46 78000.000000
Rwneg34_47 in34_47 sn34_47 202000.000000
Rwneg34_48 in34_48 sn34_48 78000.000000
Rwneg34_49 in34_49 sn34_49 202000.000000
Rwneg34_50 in34_50 sn34_50 78000.000000
Rwneg34_51 in34_51 sn34_51 202000.000000
Rwneg34_52 in34_52 sn34_52 78000.000000
Rwneg34_53 in34_53 sn34_53 78000.000000
Rwneg34_54 in34_54 sn34_54 202000.000000
Rwneg34_55 in34_55 sn34_55 78000.000000
Rwneg34_56 in34_56 sn34_56 202000.000000
Rwneg34_57 in34_57 sn34_57 202000.000000
Rwneg34_58 in34_58 sn34_58 78000.000000
Rwneg34_59 in34_59 sn34_59 202000.000000
Rwneg34_60 in34_60 sn34_60 78000.000000
Rwneg34_61 in34_61 sn34_61 78000.000000
Rwneg34_62 in34_62 sn34_62 78000.000000
Rwneg34_63 in34_63 sn34_63 202000.000000
Rwneg34_64 in34_64 sn34_64 202000.000000
Rwneg34_65 in34_65 sn34_65 202000.000000
Rwneg34_66 in34_66 sn34_66 78000.000000
Rwneg34_67 in34_67 sn34_67 202000.000000
Rwneg34_68 in34_68 sn34_68 202000.000000
Rwneg34_69 in34_69 sn34_69 202000.000000
Rwneg34_70 in34_70 sn34_70 78000.000000
Rwneg34_71 in34_71 sn34_71 202000.000000
Rwneg34_72 in34_72 sn34_72 202000.000000
Rwneg34_73 in34_73 sn34_73 78000.000000
Rwneg34_74 in34_74 sn34_74 78000.000000
Rwneg34_75 in34_75 sn34_75 202000.000000
Rwneg34_76 in34_76 sn34_76 78000.000000
Rwneg34_77 in34_77 sn34_77 202000.000000
Rwneg34_78 in34_78 sn34_78 202000.000000
Rwneg34_79 in34_79 sn34_79 202000.000000
Rwneg34_80 in34_80 sn34_80 78000.000000
Rwneg34_81 in34_81 sn34_81 78000.000000
Rwneg34_82 in34_82 sn34_82 202000.000000
Rwneg34_83 in34_83 sn34_83 78000.000000
Rwneg34_84 in34_84 sn34_84 78000.000000
Rwneg35_1 in35_1 sn35_1 202000.000000
Rwneg35_2 in35_2 sn35_2 202000.000000
Rwneg35_3 in35_3 sn35_3 202000.000000
Rwneg35_4 in35_4 sn35_4 78000.000000
Rwneg35_5 in35_5 sn35_5 202000.000000
Rwneg35_6 in35_6 sn35_6 202000.000000
Rwneg35_7 in35_7 sn35_7 202000.000000
Rwneg35_8 in35_8 sn35_8 78000.000000
Rwneg35_9 in35_9 sn35_9 202000.000000
Rwneg35_10 in35_10 sn35_10 202000.000000
Rwneg35_11 in35_11 sn35_11 202000.000000
Rwneg35_12 in35_12 sn35_12 78000.000000
Rwneg35_13 in35_13 sn35_13 78000.000000
Rwneg35_14 in35_14 sn35_14 202000.000000
Rwneg35_15 in35_15 sn35_15 202000.000000
Rwneg35_16 in35_16 sn35_16 202000.000000
Rwneg35_17 in35_17 sn35_17 202000.000000
Rwneg35_18 in35_18 sn35_18 78000.000000
Rwneg35_19 in35_19 sn35_19 202000.000000
Rwneg35_20 in35_20 sn35_20 202000.000000
Rwneg35_21 in35_21 sn35_21 202000.000000
Rwneg35_22 in35_22 sn35_22 202000.000000
Rwneg35_23 in35_23 sn35_23 78000.000000
Rwneg35_24 in35_24 sn35_24 202000.000000
Rwneg35_25 in35_25 sn35_25 78000.000000
Rwneg35_26 in35_26 sn35_26 78000.000000
Rwneg35_27 in35_27 sn35_27 78000.000000
Rwneg35_28 in35_28 sn35_28 202000.000000
Rwneg35_29 in35_29 sn35_29 202000.000000
Rwneg35_30 in35_30 sn35_30 78000.000000
Rwneg35_31 in35_31 sn35_31 78000.000000
Rwneg35_32 in35_32 sn35_32 202000.000000
Rwneg35_33 in35_33 sn35_33 202000.000000
Rwneg35_34 in35_34 sn35_34 78000.000000
Rwneg35_35 in35_35 sn35_35 78000.000000
Rwneg35_36 in35_36 sn35_36 78000.000000
Rwneg35_37 in35_37 sn35_37 202000.000000
Rwneg35_38 in35_38 sn35_38 202000.000000
Rwneg35_39 in35_39 sn35_39 78000.000000
Rwneg35_40 in35_40 sn35_40 202000.000000
Rwneg35_41 in35_41 sn35_41 202000.000000
Rwneg35_42 in35_42 sn35_42 202000.000000
Rwneg35_43 in35_43 sn35_43 202000.000000
Rwneg35_44 in35_44 sn35_44 202000.000000
Rwneg35_45 in35_45 sn35_45 202000.000000
Rwneg35_46 in35_46 sn35_46 78000.000000
Rwneg35_47 in35_47 sn35_47 202000.000000
Rwneg35_48 in35_48 sn35_48 78000.000000
Rwneg35_49 in35_49 sn35_49 202000.000000
Rwneg35_50 in35_50 sn35_50 202000.000000
Rwneg35_51 in35_51 sn35_51 202000.000000
Rwneg35_52 in35_52 sn35_52 202000.000000
Rwneg35_53 in35_53 sn35_53 78000.000000
Rwneg35_54 in35_54 sn35_54 78000.000000
Rwneg35_55 in35_55 sn35_55 78000.000000
Rwneg35_56 in35_56 sn35_56 78000.000000
Rwneg35_57 in35_57 sn35_57 202000.000000
Rwneg35_58 in35_58 sn35_58 202000.000000
Rwneg35_59 in35_59 sn35_59 78000.000000
Rwneg35_60 in35_60 sn35_60 78000.000000
Rwneg35_61 in35_61 sn35_61 78000.000000
Rwneg35_62 in35_62 sn35_62 202000.000000
Rwneg35_63 in35_63 sn35_63 78000.000000
Rwneg35_64 in35_64 sn35_64 78000.000000
Rwneg35_65 in35_65 sn35_65 78000.000000
Rwneg35_66 in35_66 sn35_66 202000.000000
Rwneg35_67 in35_67 sn35_67 78000.000000
Rwneg35_68 in35_68 sn35_68 78000.000000
Rwneg35_69 in35_69 sn35_69 78000.000000
Rwneg35_70 in35_70 sn35_70 78000.000000
Rwneg35_71 in35_71 sn35_71 78000.000000
Rwneg35_72 in35_72 sn35_72 202000.000000
Rwneg35_73 in35_73 sn35_73 78000.000000
Rwneg35_74 in35_74 sn35_74 78000.000000
Rwneg35_75 in35_75 sn35_75 202000.000000
Rwneg35_76 in35_76 sn35_76 78000.000000
Rwneg35_77 in35_77 sn35_77 78000.000000
Rwneg35_78 in35_78 sn35_78 202000.000000
Rwneg35_79 in35_79 sn35_79 78000.000000
Rwneg35_80 in35_80 sn35_80 78000.000000
Rwneg35_81 in35_81 sn35_81 78000.000000
Rwneg35_82 in35_82 sn35_82 78000.000000
Rwneg35_83 in35_83 sn35_83 78000.000000
Rwneg35_84 in35_84 sn35_84 78000.000000
Rwneg36_1 in36_1 sn36_1 202000.000000
Rwneg36_2 in36_2 sn36_2 202000.000000
Rwneg36_3 in36_3 sn36_3 202000.000000
Rwneg36_4 in36_4 sn36_4 78000.000000
Rwneg36_5 in36_5 sn36_5 78000.000000
Rwneg36_6 in36_6 sn36_6 78000.000000
Rwneg36_7 in36_7 sn36_7 202000.000000
Rwneg36_8 in36_8 sn36_8 202000.000000
Rwneg36_9 in36_9 sn36_9 78000.000000
Rwneg36_10 in36_10 sn36_10 202000.000000
Rwneg36_11 in36_11 sn36_11 78000.000000
Rwneg36_12 in36_12 sn36_12 78000.000000
Rwneg36_13 in36_13 sn36_13 78000.000000
Rwneg36_14 in36_14 sn36_14 78000.000000
Rwneg36_15 in36_15 sn36_15 78000.000000
Rwneg36_16 in36_16 sn36_16 78000.000000
Rwneg36_17 in36_17 sn36_17 78000.000000
Rwneg36_18 in36_18 sn36_18 78000.000000
Rwneg36_19 in36_19 sn36_19 78000.000000
Rwneg36_20 in36_20 sn36_20 202000.000000
Rwneg36_21 in36_21 sn36_21 78000.000000
Rwneg36_22 in36_22 sn36_22 78000.000000
Rwneg36_23 in36_23 sn36_23 202000.000000
Rwneg36_24 in36_24 sn36_24 202000.000000
Rwneg36_25 in36_25 sn36_25 202000.000000
Rwneg36_26 in36_26 sn36_26 202000.000000
Rwneg36_27 in36_27 sn36_27 78000.000000
Rwneg36_28 in36_28 sn36_28 202000.000000
Rwneg36_29 in36_29 sn36_29 202000.000000
Rwneg36_30 in36_30 sn36_30 78000.000000
Rwneg36_31 in36_31 sn36_31 78000.000000
Rwneg36_32 in36_32 sn36_32 78000.000000
Rwneg36_33 in36_33 sn36_33 202000.000000
Rwneg36_34 in36_34 sn36_34 78000.000000
Rwneg36_35 in36_35 sn36_35 202000.000000
Rwneg36_36 in36_36 sn36_36 202000.000000
Rwneg36_37 in36_37 sn36_37 202000.000000
Rwneg36_38 in36_38 sn36_38 78000.000000
Rwneg36_39 in36_39 sn36_39 78000.000000
Rwneg36_40 in36_40 sn36_40 78000.000000
Rwneg36_41 in36_41 sn36_41 78000.000000
Rwneg36_42 in36_42 sn36_42 202000.000000
Rwneg36_43 in36_43 sn36_43 202000.000000
Rwneg36_44 in36_44 sn36_44 202000.000000
Rwneg36_45 in36_45 sn36_45 78000.000000
Rwneg36_46 in36_46 sn36_46 202000.000000
Rwneg36_47 in36_47 sn36_47 202000.000000
Rwneg36_48 in36_48 sn36_48 202000.000000
Rwneg36_49 in36_49 sn36_49 202000.000000
Rwneg36_50 in36_50 sn36_50 202000.000000
Rwneg36_51 in36_51 sn36_51 202000.000000
Rwneg36_52 in36_52 sn36_52 202000.000000
Rwneg36_53 in36_53 sn36_53 202000.000000
Rwneg36_54 in36_54 sn36_54 78000.000000
Rwneg36_55 in36_55 sn36_55 78000.000000
Rwneg36_56 in36_56 sn36_56 202000.000000
Rwneg36_57 in36_57 sn36_57 78000.000000
Rwneg36_58 in36_58 sn36_58 78000.000000
Rwneg36_59 in36_59 sn36_59 78000.000000
Rwneg36_60 in36_60 sn36_60 202000.000000
Rwneg36_61 in36_61 sn36_61 202000.000000
Rwneg36_62 in36_62 sn36_62 202000.000000
Rwneg36_63 in36_63 sn36_63 202000.000000
Rwneg36_64 in36_64 sn36_64 78000.000000
Rwneg36_65 in36_65 sn36_65 202000.000000
Rwneg36_66 in36_66 sn36_66 202000.000000
Rwneg36_67 in36_67 sn36_67 78000.000000
Rwneg36_68 in36_68 sn36_68 78000.000000
Rwneg36_69 in36_69 sn36_69 202000.000000
Rwneg36_70 in36_70 sn36_70 202000.000000
Rwneg36_71 in36_71 sn36_71 202000.000000
Rwneg36_72 in36_72 sn36_72 202000.000000
Rwneg36_73 in36_73 sn36_73 78000.000000
Rwneg36_74 in36_74 sn36_74 78000.000000
Rwneg36_75 in36_75 sn36_75 78000.000000
Rwneg36_76 in36_76 sn36_76 202000.000000
Rwneg36_77 in36_77 sn36_77 78000.000000
Rwneg36_78 in36_78 sn36_78 202000.000000
Rwneg36_79 in36_79 sn36_79 202000.000000
Rwneg36_80 in36_80 sn36_80 78000.000000
Rwneg36_81 in36_81 sn36_81 202000.000000
Rwneg36_82 in36_82 sn36_82 202000.000000
Rwneg36_83 in36_83 sn36_83 78000.000000
Rwneg36_84 in36_84 sn36_84 78000.000000
Rwneg37_1 in37_1 sn37_1 202000.000000
Rwneg37_2 in37_2 sn37_2 78000.000000
Rwneg37_3 in37_3 sn37_3 202000.000000
Rwneg37_4 in37_4 sn37_4 78000.000000
Rwneg37_5 in37_5 sn37_5 202000.000000
Rwneg37_6 in37_6 sn37_6 202000.000000
Rwneg37_7 in37_7 sn37_7 78000.000000
Rwneg37_8 in37_8 sn37_8 78000.000000
Rwneg37_9 in37_9 sn37_9 202000.000000
Rwneg37_10 in37_10 sn37_10 202000.000000
Rwneg37_11 in37_11 sn37_11 78000.000000
Rwneg37_12 in37_12 sn37_12 202000.000000
Rwneg37_13 in37_13 sn37_13 202000.000000
Rwneg37_14 in37_14 sn37_14 202000.000000
Rwneg37_15 in37_15 sn37_15 202000.000000
Rwneg37_16 in37_16 sn37_16 202000.000000
Rwneg37_17 in37_17 sn37_17 78000.000000
Rwneg37_18 in37_18 sn37_18 202000.000000
Rwneg37_19 in37_19 sn37_19 202000.000000
Rwneg37_20 in37_20 sn37_20 202000.000000
Rwneg37_21 in37_21 sn37_21 202000.000000
Rwneg37_22 in37_22 sn37_22 202000.000000
Rwneg37_23 in37_23 sn37_23 78000.000000
Rwneg37_24 in37_24 sn37_24 202000.000000
Rwneg37_25 in37_25 sn37_25 78000.000000
Rwneg37_26 in37_26 sn37_26 78000.000000
Rwneg37_27 in37_27 sn37_27 202000.000000
Rwneg37_28 in37_28 sn37_28 202000.000000
Rwneg37_29 in37_29 sn37_29 202000.000000
Rwneg37_30 in37_30 sn37_30 202000.000000
Rwneg37_31 in37_31 sn37_31 202000.000000
Rwneg37_32 in37_32 sn37_32 78000.000000
Rwneg37_33 in37_33 sn37_33 78000.000000
Rwneg37_34 in37_34 sn37_34 202000.000000
Rwneg37_35 in37_35 sn37_35 202000.000000
Rwneg37_36 in37_36 sn37_36 202000.000000
Rwneg37_37 in37_37 sn37_37 78000.000000
Rwneg37_38 in37_38 sn37_38 202000.000000
Rwneg37_39 in37_39 sn37_39 202000.000000
Rwneg37_40 in37_40 sn37_40 202000.000000
Rwneg37_41 in37_41 sn37_41 78000.000000
Rwneg37_42 in37_42 sn37_42 78000.000000
Rwneg37_43 in37_43 sn37_43 78000.000000
Rwneg37_44 in37_44 sn37_44 78000.000000
Rwneg37_45 in37_45 sn37_45 202000.000000
Rwneg37_46 in37_46 sn37_46 202000.000000
Rwneg37_47 in37_47 sn37_47 202000.000000
Rwneg37_48 in37_48 sn37_48 202000.000000
Rwneg37_49 in37_49 sn37_49 202000.000000
Rwneg37_50 in37_50 sn37_50 202000.000000
Rwneg37_51 in37_51 sn37_51 78000.000000
Rwneg37_52 in37_52 sn37_52 202000.000000
Rwneg37_53 in37_53 sn37_53 78000.000000
Rwneg37_54 in37_54 sn37_54 78000.000000
Rwneg37_55 in37_55 sn37_55 78000.000000
Rwneg37_56 in37_56 sn37_56 78000.000000
Rwneg37_57 in37_57 sn37_57 202000.000000
Rwneg37_58 in37_58 sn37_58 78000.000000
Rwneg37_59 in37_59 sn37_59 202000.000000
Rwneg37_60 in37_60 sn37_60 78000.000000
Rwneg37_61 in37_61 sn37_61 202000.000000
Rwneg37_62 in37_62 sn37_62 78000.000000
Rwneg37_63 in37_63 sn37_63 78000.000000
Rwneg37_64 in37_64 sn37_64 78000.000000
Rwneg37_65 in37_65 sn37_65 202000.000000
Rwneg37_66 in37_66 sn37_66 78000.000000
Rwneg37_67 in37_67 sn37_67 202000.000000
Rwneg37_68 in37_68 sn37_68 78000.000000
Rwneg37_69 in37_69 sn37_69 78000.000000
Rwneg37_70 in37_70 sn37_70 202000.000000
Rwneg37_71 in37_71 sn37_71 78000.000000
Rwneg37_72 in37_72 sn37_72 202000.000000
Rwneg37_73 in37_73 sn37_73 202000.000000
Rwneg37_74 in37_74 sn37_74 202000.000000
Rwneg37_75 in37_75 sn37_75 202000.000000
Rwneg37_76 in37_76 sn37_76 202000.000000
Rwneg37_77 in37_77 sn37_77 202000.000000
Rwneg37_78 in37_78 sn37_78 202000.000000
Rwneg37_79 in37_79 sn37_79 78000.000000
Rwneg37_80 in37_80 sn37_80 78000.000000
Rwneg37_81 in37_81 sn37_81 78000.000000
Rwneg37_82 in37_82 sn37_82 78000.000000
Rwneg37_83 in37_83 sn37_83 78000.000000
Rwneg37_84 in37_84 sn37_84 78000.000000
Rwneg38_1 in38_1 sn38_1 202000.000000
Rwneg38_2 in38_2 sn38_2 78000.000000
Rwneg38_3 in38_3 sn38_3 78000.000000
Rwneg38_4 in38_4 sn38_4 78000.000000
Rwneg38_5 in38_5 sn38_5 78000.000000
Rwneg38_6 in38_6 sn38_6 202000.000000
Rwneg38_7 in38_7 sn38_7 78000.000000
Rwneg38_8 in38_8 sn38_8 78000.000000
Rwneg38_9 in38_9 sn38_9 78000.000000
Rwneg38_10 in38_10 sn38_10 78000.000000
Rwneg38_11 in38_11 sn38_11 202000.000000
Rwneg38_12 in38_12 sn38_12 78000.000000
Rwneg38_13 in38_13 sn38_13 202000.000000
Rwneg38_14 in38_14 sn38_14 78000.000000
Rwneg38_15 in38_15 sn38_15 202000.000000
Rwneg38_16 in38_16 sn38_16 78000.000000
Rwneg38_17 in38_17 sn38_17 202000.000000
Rwneg38_18 in38_18 sn38_18 78000.000000
Rwneg38_19 in38_19 sn38_19 78000.000000
Rwneg38_20 in38_20 sn38_20 202000.000000
Rwneg38_21 in38_21 sn38_21 202000.000000
Rwneg38_22 in38_22 sn38_22 202000.000000
Rwneg38_23 in38_23 sn38_23 202000.000000
Rwneg38_24 in38_24 sn38_24 202000.000000
Rwneg38_25 in38_25 sn38_25 202000.000000
Rwneg38_26 in38_26 sn38_26 202000.000000
Rwneg38_27 in38_27 sn38_27 78000.000000
Rwneg38_28 in38_28 sn38_28 78000.000000
Rwneg38_29 in38_29 sn38_29 78000.000000
Rwneg38_30 in38_30 sn38_30 78000.000000
Rwneg38_31 in38_31 sn38_31 202000.000000
Rwneg38_32 in38_32 sn38_32 202000.000000
Rwneg38_33 in38_33 sn38_33 202000.000000
Rwneg38_34 in38_34 sn38_34 78000.000000
Rwneg38_35 in38_35 sn38_35 78000.000000
Rwneg38_36 in38_36 sn38_36 78000.000000
Rwneg38_37 in38_37 sn38_37 202000.000000
Rwneg38_38 in38_38 sn38_38 78000.000000
Rwneg38_39 in38_39 sn38_39 78000.000000
Rwneg38_40 in38_40 sn38_40 202000.000000
Rwneg38_41 in38_41 sn38_41 78000.000000
Rwneg38_42 in38_42 sn38_42 202000.000000
Rwneg38_43 in38_43 sn38_43 202000.000000
Rwneg38_44 in38_44 sn38_44 202000.000000
Rwneg38_45 in38_45 sn38_45 78000.000000
Rwneg38_46 in38_46 sn38_46 78000.000000
Rwneg38_47 in38_47 sn38_47 78000.000000
Rwneg38_48 in38_48 sn38_48 78000.000000
Rwneg38_49 in38_49 sn38_49 78000.000000
Rwneg38_50 in38_50 sn38_50 78000.000000
Rwneg38_51 in38_51 sn38_51 202000.000000
Rwneg38_52 in38_52 sn38_52 78000.000000
Rwneg38_53 in38_53 sn38_53 78000.000000
Rwneg38_54 in38_54 sn38_54 202000.000000
Rwneg38_55 in38_55 sn38_55 78000.000000
Rwneg38_56 in38_56 sn38_56 202000.000000
Rwneg38_57 in38_57 sn38_57 202000.000000
Rwneg38_58 in38_58 sn38_58 202000.000000
Rwneg38_59 in38_59 sn38_59 78000.000000
Rwneg38_60 in38_60 sn38_60 78000.000000
Rwneg38_61 in38_61 sn38_61 78000.000000
Rwneg38_62 in38_62 sn38_62 202000.000000
Rwneg38_63 in38_63 sn38_63 78000.000000
Rwneg38_64 in38_64 sn38_64 202000.000000
Rwneg38_65 in38_65 sn38_65 78000.000000
Rwneg38_66 in38_66 sn38_66 78000.000000
Rwneg38_67 in38_67 sn38_67 78000.000000
Rwneg38_68 in38_68 sn38_68 202000.000000
Rwneg38_69 in38_69 sn38_69 78000.000000
Rwneg38_70 in38_70 sn38_70 202000.000000
Rwneg38_71 in38_71 sn38_71 78000.000000
Rwneg38_72 in38_72 sn38_72 202000.000000
Rwneg38_73 in38_73 sn38_73 202000.000000
Rwneg38_74 in38_74 sn38_74 78000.000000
Rwneg38_75 in38_75 sn38_75 78000.000000
Rwneg38_76 in38_76 sn38_76 78000.000000
Rwneg38_77 in38_77 sn38_77 78000.000000
Rwneg38_78 in38_78 sn38_78 78000.000000
Rwneg38_79 in38_79 sn38_79 78000.000000
Rwneg38_80 in38_80 sn38_80 202000.000000
Rwneg38_81 in38_81 sn38_81 202000.000000
Rwneg38_82 in38_82 sn38_82 78000.000000
Rwneg38_83 in38_83 sn38_83 78000.000000
Rwneg38_84 in38_84 sn38_84 78000.000000
Rwneg39_1 in39_1 sn39_1 202000.000000
Rwneg39_2 in39_2 sn39_2 202000.000000
Rwneg39_3 in39_3 sn39_3 202000.000000
Rwneg39_4 in39_4 sn39_4 202000.000000
Rwneg39_5 in39_5 sn39_5 202000.000000
Rwneg39_6 in39_6 sn39_6 202000.000000
Rwneg39_7 in39_7 sn39_7 78000.000000
Rwneg39_8 in39_8 sn39_8 202000.000000
Rwneg39_9 in39_9 sn39_9 202000.000000
Rwneg39_10 in39_10 sn39_10 78000.000000
Rwneg39_11 in39_11 sn39_11 78000.000000
Rwneg39_12 in39_12 sn39_12 78000.000000
Rwneg39_13 in39_13 sn39_13 202000.000000
Rwneg39_14 in39_14 sn39_14 202000.000000
Rwneg39_15 in39_15 sn39_15 78000.000000
Rwneg39_16 in39_16 sn39_16 202000.000000
Rwneg39_17 in39_17 sn39_17 78000.000000
Rwneg39_18 in39_18 sn39_18 202000.000000
Rwneg39_19 in39_19 sn39_19 78000.000000
Rwneg39_20 in39_20 sn39_20 202000.000000
Rwneg39_21 in39_21 sn39_21 78000.000000
Rwneg39_22 in39_22 sn39_22 78000.000000
Rwneg39_23 in39_23 sn39_23 202000.000000
Rwneg39_24 in39_24 sn39_24 78000.000000
Rwneg39_25 in39_25 sn39_25 202000.000000
Rwneg39_26 in39_26 sn39_26 202000.000000
Rwneg39_27 in39_27 sn39_27 202000.000000
Rwneg39_28 in39_28 sn39_28 78000.000000
Rwneg39_29 in39_29 sn39_29 202000.000000
Rwneg39_30 in39_30 sn39_30 202000.000000
Rwneg39_31 in39_31 sn39_31 78000.000000
Rwneg39_32 in39_32 sn39_32 202000.000000
Rwneg39_33 in39_33 sn39_33 78000.000000
Rwneg39_34 in39_34 sn39_34 78000.000000
Rwneg39_35 in39_35 sn39_35 202000.000000
Rwneg39_36 in39_36 sn39_36 78000.000000
Rwneg39_37 in39_37 sn39_37 78000.000000
Rwneg39_38 in39_38 sn39_38 78000.000000
Rwneg39_39 in39_39 sn39_39 202000.000000
Rwneg39_40 in39_40 sn39_40 78000.000000
Rwneg39_41 in39_41 sn39_41 202000.000000
Rwneg39_42 in39_42 sn39_42 202000.000000
Rwneg39_43 in39_43 sn39_43 78000.000000
Rwneg39_44 in39_44 sn39_44 202000.000000
Rwneg39_45 in39_45 sn39_45 202000.000000
Rwneg39_46 in39_46 sn39_46 202000.000000
Rwneg39_47 in39_47 sn39_47 202000.000000
Rwneg39_48 in39_48 sn39_48 78000.000000
Rwneg39_49 in39_49 sn39_49 78000.000000
Rwneg39_50 in39_50 sn39_50 78000.000000
Rwneg39_51 in39_51 sn39_51 78000.000000
Rwneg39_52 in39_52 sn39_52 78000.000000
Rwneg39_53 in39_53 sn39_53 202000.000000
Rwneg39_54 in39_54 sn39_54 202000.000000
Rwneg39_55 in39_55 sn39_55 78000.000000
Rwneg39_56 in39_56 sn39_56 202000.000000
Rwneg39_57 in39_57 sn39_57 78000.000000
Rwneg39_58 in39_58 sn39_58 202000.000000
Rwneg39_59 in39_59 sn39_59 202000.000000
Rwneg39_60 in39_60 sn39_60 202000.000000
Rwneg39_61 in39_61 sn39_61 78000.000000
Rwneg39_62 in39_62 sn39_62 78000.000000
Rwneg39_63 in39_63 sn39_63 78000.000000
Rwneg39_64 in39_64 sn39_64 78000.000000
Rwneg39_65 in39_65 sn39_65 78000.000000
Rwneg39_66 in39_66 sn39_66 202000.000000
Rwneg39_67 in39_67 sn39_67 78000.000000
Rwneg39_68 in39_68 sn39_68 78000.000000
Rwneg39_69 in39_69 sn39_69 78000.000000
Rwneg39_70 in39_70 sn39_70 78000.000000
Rwneg39_71 in39_71 sn39_71 202000.000000
Rwneg39_72 in39_72 sn39_72 202000.000000
Rwneg39_73 in39_73 sn39_73 78000.000000
Rwneg39_74 in39_74 sn39_74 202000.000000
Rwneg39_75 in39_75 sn39_75 202000.000000
Rwneg39_76 in39_76 sn39_76 202000.000000
Rwneg39_77 in39_77 sn39_77 202000.000000
Rwneg39_78 in39_78 sn39_78 202000.000000
Rwneg39_79 in39_79 sn39_79 202000.000000
Rwneg39_80 in39_80 sn39_80 202000.000000
Rwneg39_81 in39_81 sn39_81 202000.000000
Rwneg39_82 in39_82 sn39_82 78000.000000
Rwneg39_83 in39_83 sn39_83 202000.000000
Rwneg39_84 in39_84 sn39_84 202000.000000
Rwneg40_1 in40_1 sn40_1 202000.000000
Rwneg40_2 in40_2 sn40_2 78000.000000
Rwneg40_3 in40_3 sn40_3 78000.000000
Rwneg40_4 in40_4 sn40_4 78000.000000
Rwneg40_5 in40_5 sn40_5 78000.000000
Rwneg40_6 in40_6 sn40_6 78000.000000
Rwneg40_7 in40_7 sn40_7 202000.000000
Rwneg40_8 in40_8 sn40_8 78000.000000
Rwneg40_9 in40_9 sn40_9 78000.000000
Rwneg40_10 in40_10 sn40_10 78000.000000
Rwneg40_11 in40_11 sn40_11 202000.000000
Rwneg40_12 in40_12 sn40_12 78000.000000
Rwneg40_13 in40_13 sn40_13 202000.000000
Rwneg40_14 in40_14 sn40_14 78000.000000
Rwneg40_15 in40_15 sn40_15 78000.000000
Rwneg40_16 in40_16 sn40_16 202000.000000
Rwneg40_17 in40_17 sn40_17 202000.000000
Rwneg40_18 in40_18 sn40_18 78000.000000
Rwneg40_19 in40_19 sn40_19 202000.000000
Rwneg40_20 in40_20 sn40_20 202000.000000
Rwneg40_21 in40_21 sn40_21 202000.000000
Rwneg40_22 in40_22 sn40_22 202000.000000
Rwneg40_23 in40_23 sn40_23 78000.000000
Rwneg40_24 in40_24 sn40_24 202000.000000
Rwneg40_25 in40_25 sn40_25 202000.000000
Rwneg40_26 in40_26 sn40_26 202000.000000
Rwneg40_27 in40_27 sn40_27 78000.000000
Rwneg40_28 in40_28 sn40_28 202000.000000
Rwneg40_29 in40_29 sn40_29 202000.000000
Rwneg40_30 in40_30 sn40_30 202000.000000
Rwneg40_31 in40_31 sn40_31 78000.000000
Rwneg40_32 in40_32 sn40_32 202000.000000
Rwneg40_33 in40_33 sn40_33 202000.000000
Rwneg40_34 in40_34 sn40_34 78000.000000
Rwneg40_35 in40_35 sn40_35 78000.000000
Rwneg40_36 in40_36 sn40_36 202000.000000
Rwneg40_37 in40_37 sn40_37 202000.000000
Rwneg40_38 in40_38 sn40_38 78000.000000
Rwneg40_39 in40_39 sn40_39 202000.000000
Rwneg40_40 in40_40 sn40_40 202000.000000
Rwneg40_41 in40_41 sn40_41 202000.000000
Rwneg40_42 in40_42 sn40_42 78000.000000
Rwneg40_43 in40_43 sn40_43 202000.000000
Rwneg40_44 in40_44 sn40_44 202000.000000
Rwneg40_45 in40_45 sn40_45 78000.000000
Rwneg40_46 in40_46 sn40_46 78000.000000
Rwneg40_47 in40_47 sn40_47 202000.000000
Rwneg40_48 in40_48 sn40_48 202000.000000
Rwneg40_49 in40_49 sn40_49 78000.000000
Rwneg40_50 in40_50 sn40_50 202000.000000
Rwneg40_51 in40_51 sn40_51 202000.000000
Rwneg40_52 in40_52 sn40_52 78000.000000
Rwneg40_53 in40_53 sn40_53 78000.000000
Rwneg40_54 in40_54 sn40_54 78000.000000
Rwneg40_55 in40_55 sn40_55 202000.000000
Rwneg40_56 in40_56 sn40_56 78000.000000
Rwneg40_57 in40_57 sn40_57 202000.000000
Rwneg40_58 in40_58 sn40_58 78000.000000
Rwneg40_59 in40_59 sn40_59 202000.000000
Rwneg40_60 in40_60 sn40_60 202000.000000
Rwneg40_61 in40_61 sn40_61 202000.000000
Rwneg40_62 in40_62 sn40_62 202000.000000
Rwneg40_63 in40_63 sn40_63 202000.000000
Rwneg40_64 in40_64 sn40_64 78000.000000
Rwneg40_65 in40_65 sn40_65 78000.000000
Rwneg40_66 in40_66 sn40_66 202000.000000
Rwneg40_67 in40_67 sn40_67 202000.000000
Rwneg40_68 in40_68 sn40_68 202000.000000
Rwneg40_69 in40_69 sn40_69 78000.000000
Rwneg40_70 in40_70 sn40_70 202000.000000
Rwneg40_71 in40_71 sn40_71 202000.000000
Rwneg40_72 in40_72 sn40_72 78000.000000
Rwneg40_73 in40_73 sn40_73 78000.000000
Rwneg40_74 in40_74 sn40_74 78000.000000
Rwneg40_75 in40_75 sn40_75 202000.000000
Rwneg40_76 in40_76 sn40_76 202000.000000
Rwneg40_77 in40_77 sn40_77 78000.000000
Rwneg40_78 in40_78 sn40_78 202000.000000
Rwneg40_79 in40_79 sn40_79 202000.000000
Rwneg40_80 in40_80 sn40_80 78000.000000
Rwneg40_81 in40_81 sn40_81 202000.000000
Rwneg40_82 in40_82 sn40_82 78000.000000
Rwneg40_83 in40_83 sn40_83 78000.000000
Rwneg40_84 in40_84 sn40_84 78000.000000
Rwneg41_1 in41_1 sn41_1 202000.000000
Rwneg41_2 in41_2 sn41_2 78000.000000
Rwneg41_3 in41_3 sn41_3 78000.000000
Rwneg41_4 in41_4 sn41_4 202000.000000
Rwneg41_5 in41_5 sn41_5 78000.000000
Rwneg41_6 in41_6 sn41_6 202000.000000
Rwneg41_7 in41_7 sn41_7 78000.000000
Rwneg41_8 in41_8 sn41_8 202000.000000
Rwneg41_9 in41_9 sn41_9 202000.000000
Rwneg41_10 in41_10 sn41_10 202000.000000
Rwneg41_11 in41_11 sn41_11 202000.000000
Rwneg41_12 in41_12 sn41_12 78000.000000
Rwneg41_13 in41_13 sn41_13 202000.000000
Rwneg41_14 in41_14 sn41_14 78000.000000
Rwneg41_15 in41_15 sn41_15 78000.000000
Rwneg41_16 in41_16 sn41_16 78000.000000
Rwneg41_17 in41_17 sn41_17 202000.000000
Rwneg41_18 in41_18 sn41_18 202000.000000
Rwneg41_19 in41_19 sn41_19 78000.000000
Rwneg41_20 in41_20 sn41_20 202000.000000
Rwneg41_21 in41_21 sn41_21 202000.000000
Rwneg41_22 in41_22 sn41_22 202000.000000
Rwneg41_23 in41_23 sn41_23 202000.000000
Rwneg41_24 in41_24 sn41_24 202000.000000
Rwneg41_25 in41_25 sn41_25 202000.000000
Rwneg41_26 in41_26 sn41_26 202000.000000
Rwneg41_27 in41_27 sn41_27 78000.000000
Rwneg41_28 in41_28 sn41_28 78000.000000
Rwneg41_29 in41_29 sn41_29 78000.000000
Rwneg41_30 in41_30 sn41_30 78000.000000
Rwneg41_31 in41_31 sn41_31 78000.000000
Rwneg41_32 in41_32 sn41_32 78000.000000
Rwneg41_33 in41_33 sn41_33 78000.000000
Rwneg41_34 in41_34 sn41_34 202000.000000
Rwneg41_35 in41_35 sn41_35 78000.000000
Rwneg41_36 in41_36 sn41_36 202000.000000
Rwneg41_37 in41_37 sn41_37 78000.000000
Rwneg41_38 in41_38 sn41_38 78000.000000
Rwneg41_39 in41_39 sn41_39 202000.000000
Rwneg41_40 in41_40 sn41_40 202000.000000
Rwneg41_41 in41_41 sn41_41 202000.000000
Rwneg41_42 in41_42 sn41_42 202000.000000
Rwneg41_43 in41_43 sn41_43 202000.000000
Rwneg41_44 in41_44 sn41_44 202000.000000
Rwneg41_45 in41_45 sn41_45 202000.000000
Rwneg41_46 in41_46 sn41_46 202000.000000
Rwneg41_47 in41_47 sn41_47 202000.000000
Rwneg41_48 in41_48 sn41_48 78000.000000
Rwneg41_49 in41_49 sn41_49 78000.000000
Rwneg41_50 in41_50 sn41_50 78000.000000
Rwneg41_51 in41_51 sn41_51 78000.000000
Rwneg41_52 in41_52 sn41_52 78000.000000
Rwneg41_53 in41_53 sn41_53 78000.000000
Rwneg41_54 in41_54 sn41_54 78000.000000
Rwneg41_55 in41_55 sn41_55 78000.000000
Rwneg41_56 in41_56 sn41_56 202000.000000
Rwneg41_57 in41_57 sn41_57 202000.000000
Rwneg41_58 in41_58 sn41_58 202000.000000
Rwneg41_59 in41_59 sn41_59 202000.000000
Rwneg41_60 in41_60 sn41_60 202000.000000
Rwneg41_61 in41_61 sn41_61 78000.000000
Rwneg41_62 in41_62 sn41_62 202000.000000
Rwneg41_63 in41_63 sn41_63 78000.000000
Rwneg41_64 in41_64 sn41_64 202000.000000
Rwneg41_65 in41_65 sn41_65 202000.000000
Rwneg41_66 in41_66 sn41_66 78000.000000
Rwneg41_67 in41_67 sn41_67 202000.000000
Rwneg41_68 in41_68 sn41_68 202000.000000
Rwneg41_69 in41_69 sn41_69 78000.000000
Rwneg41_70 in41_70 sn41_70 202000.000000
Rwneg41_71 in41_71 sn41_71 202000.000000
Rwneg41_72 in41_72 sn41_72 78000.000000
Rwneg41_73 in41_73 sn41_73 78000.000000
Rwneg41_74 in41_74 sn41_74 78000.000000
Rwneg41_75 in41_75 sn41_75 202000.000000
Rwneg41_76 in41_76 sn41_76 78000.000000
Rwneg41_77 in41_77 sn41_77 202000.000000
Rwneg41_78 in41_78 sn41_78 78000.000000
Rwneg41_79 in41_79 sn41_79 78000.000000
Rwneg41_80 in41_80 sn41_80 202000.000000
Rwneg41_81 in41_81 sn41_81 202000.000000
Rwneg41_82 in41_82 sn41_82 78000.000000
Rwneg41_83 in41_83 sn41_83 202000.000000
Rwneg41_84 in41_84 sn41_84 202000.000000
Rwneg42_1 in42_1 sn42_1 202000.000000
Rwneg42_2 in42_2 sn42_2 78000.000000
Rwneg42_3 in42_3 sn42_3 202000.000000
Rwneg42_4 in42_4 sn42_4 202000.000000
Rwneg42_5 in42_5 sn42_5 202000.000000
Rwneg42_6 in42_6 sn42_6 202000.000000
Rwneg42_7 in42_7 sn42_7 202000.000000
Rwneg42_8 in42_8 sn42_8 202000.000000
Rwneg42_9 in42_9 sn42_9 202000.000000
Rwneg42_10 in42_10 sn42_10 202000.000000
Rwneg42_11 in42_11 sn42_11 78000.000000
Rwneg42_12 in42_12 sn42_12 202000.000000
Rwneg42_13 in42_13 sn42_13 202000.000000
Rwneg42_14 in42_14 sn42_14 78000.000000
Rwneg42_15 in42_15 sn42_15 202000.000000
Rwneg42_16 in42_16 sn42_16 202000.000000
Rwneg42_17 in42_17 sn42_17 78000.000000
Rwneg42_18 in42_18 sn42_18 202000.000000
Rwneg42_19 in42_19 sn42_19 202000.000000
Rwneg42_20 in42_20 sn42_20 202000.000000
Rwneg42_21 in42_21 sn42_21 78000.000000
Rwneg42_22 in42_22 sn42_22 202000.000000
Rwneg42_23 in42_23 sn42_23 78000.000000
Rwneg42_24 in42_24 sn42_24 78000.000000
Rwneg42_25 in42_25 sn42_25 202000.000000
Rwneg42_26 in42_26 sn42_26 202000.000000
Rwneg42_27 in42_27 sn42_27 202000.000000
Rwneg42_28 in42_28 sn42_28 202000.000000
Rwneg42_29 in42_29 sn42_29 78000.000000
Rwneg42_30 in42_30 sn42_30 202000.000000
Rwneg42_31 in42_31 sn42_31 78000.000000
Rwneg42_32 in42_32 sn42_32 78000.000000
Rwneg42_33 in42_33 sn42_33 202000.000000
Rwneg42_34 in42_34 sn42_34 202000.000000
Rwneg42_35 in42_35 sn42_35 202000.000000
Rwneg42_36 in42_36 sn42_36 202000.000000
Rwneg42_37 in42_37 sn42_37 78000.000000
Rwneg42_38 in42_38 sn42_38 202000.000000
Rwneg42_39 in42_39 sn42_39 202000.000000
Rwneg42_40 in42_40 sn42_40 78000.000000
Rwneg42_41 in42_41 sn42_41 78000.000000
Rwneg42_42 in42_42 sn42_42 78000.000000
Rwneg42_43 in42_43 sn42_43 202000.000000
Rwneg42_44 in42_44 sn42_44 78000.000000
Rwneg42_45 in42_45 sn42_45 202000.000000
Rwneg42_46 in42_46 sn42_46 78000.000000
Rwneg42_47 in42_47 sn42_47 202000.000000
Rwneg42_48 in42_48 sn42_48 78000.000000
Rwneg42_49 in42_49 sn42_49 78000.000000
Rwneg42_50 in42_50 sn42_50 78000.000000
Rwneg42_51 in42_51 sn42_51 78000.000000
Rwneg42_52 in42_52 sn42_52 78000.000000
Rwneg42_53 in42_53 sn42_53 202000.000000
Rwneg42_54 in42_54 sn42_54 202000.000000
Rwneg42_55 in42_55 sn42_55 78000.000000
Rwneg42_56 in42_56 sn42_56 202000.000000
Rwneg42_57 in42_57 sn42_57 202000.000000
Rwneg42_58 in42_58 sn42_58 78000.000000
Rwneg42_59 in42_59 sn42_59 78000.000000
Rwneg42_60 in42_60 sn42_60 202000.000000
Rwneg42_61 in42_61 sn42_61 78000.000000
Rwneg42_62 in42_62 sn42_62 78000.000000
Rwneg42_63 in42_63 sn42_63 202000.000000
Rwneg42_64 in42_64 sn42_64 78000.000000
Rwneg42_65 in42_65 sn42_65 202000.000000
Rwneg42_66 in42_66 sn42_66 78000.000000
Rwneg42_67 in42_67 sn42_67 78000.000000
Rwneg42_68 in42_68 sn42_68 78000.000000
Rwneg42_69 in42_69 sn42_69 78000.000000
Rwneg42_70 in42_70 sn42_70 78000.000000
Rwneg42_71 in42_71 sn42_71 202000.000000
Rwneg42_72 in42_72 sn42_72 202000.000000
Rwneg42_73 in42_73 sn42_73 78000.000000
Rwneg42_74 in42_74 sn42_74 78000.000000
Rwneg42_75 in42_75 sn42_75 202000.000000
Rwneg42_76 in42_76 sn42_76 78000.000000
Rwneg42_77 in42_77 sn42_77 202000.000000
Rwneg42_78 in42_78 sn42_78 78000.000000
Rwneg42_79 in42_79 sn42_79 78000.000000
Rwneg42_80 in42_80 sn42_80 202000.000000
Rwneg42_81 in42_81 sn42_81 78000.000000
Rwneg42_82 in42_82 sn42_82 202000.000000
Rwneg42_83 in42_83 sn42_83 202000.000000
Rwneg42_84 in42_84 sn42_84 202000.000000
Rwneg43_1 in43_1 sn43_1 202000.000000
Rwneg43_2 in43_2 sn43_2 78000.000000
Rwneg43_3 in43_3 sn43_3 78000.000000
Rwneg43_4 in43_4 sn43_4 202000.000000
Rwneg43_5 in43_5 sn43_5 202000.000000
Rwneg43_6 in43_6 sn43_6 78000.000000
Rwneg43_7 in43_7 sn43_7 202000.000000
Rwneg43_8 in43_8 sn43_8 202000.000000
Rwneg43_9 in43_9 sn43_9 202000.000000
Rwneg43_10 in43_10 sn43_10 202000.000000
Rwneg43_11 in43_11 sn43_11 78000.000000
Rwneg43_12 in43_12 sn43_12 78000.000000
Rwneg43_13 in43_13 sn43_13 202000.000000
Rwneg43_14 in43_14 sn43_14 202000.000000
Rwneg43_15 in43_15 sn43_15 78000.000000
Rwneg43_16 in43_16 sn43_16 202000.000000
Rwneg43_17 in43_17 sn43_17 78000.000000
Rwneg43_18 in43_18 sn43_18 78000.000000
Rwneg43_19 in43_19 sn43_19 202000.000000
Rwneg43_20 in43_20 sn43_20 202000.000000
Rwneg43_21 in43_21 sn43_21 78000.000000
Rwneg43_22 in43_22 sn43_22 202000.000000
Rwneg43_23 in43_23 sn43_23 78000.000000
Rwneg43_24 in43_24 sn43_24 78000.000000
Rwneg43_25 in43_25 sn43_25 78000.000000
Rwneg43_26 in43_26 sn43_26 202000.000000
Rwneg43_27 in43_27 sn43_27 202000.000000
Rwneg43_28 in43_28 sn43_28 202000.000000
Rwneg43_29 in43_29 sn43_29 202000.000000
Rwneg43_30 in43_30 sn43_30 78000.000000
Rwneg43_31 in43_31 sn43_31 202000.000000
Rwneg43_32 in43_32 sn43_32 202000.000000
Rwneg43_33 in43_33 sn43_33 78000.000000
Rwneg43_34 in43_34 sn43_34 202000.000000
Rwneg43_35 in43_35 sn43_35 78000.000000
Rwneg43_36 in43_36 sn43_36 202000.000000
Rwneg43_37 in43_37 sn43_37 202000.000000
Rwneg43_38 in43_38 sn43_38 202000.000000
Rwneg43_39 in43_39 sn43_39 202000.000000
Rwneg43_40 in43_40 sn43_40 202000.000000
Rwneg43_41 in43_41 sn43_41 202000.000000
Rwneg43_42 in43_42 sn43_42 78000.000000
Rwneg43_43 in43_43 sn43_43 78000.000000
Rwneg43_44 in43_44 sn43_44 78000.000000
Rwneg43_45 in43_45 sn43_45 202000.000000
Rwneg43_46 in43_46 sn43_46 202000.000000
Rwneg43_47 in43_47 sn43_47 78000.000000
Rwneg43_48 in43_48 sn43_48 78000.000000
Rwneg43_49 in43_49 sn43_49 202000.000000
Rwneg43_50 in43_50 sn43_50 202000.000000
Rwneg43_51 in43_51 sn43_51 78000.000000
Rwneg43_52 in43_52 sn43_52 202000.000000
Rwneg43_53 in43_53 sn43_53 202000.000000
Rwneg43_54 in43_54 sn43_54 202000.000000
Rwneg43_55 in43_55 sn43_55 202000.000000
Rwneg43_56 in43_56 sn43_56 202000.000000
Rwneg43_57 in43_57 sn43_57 78000.000000
Rwneg43_58 in43_58 sn43_58 202000.000000
Rwneg43_59 in43_59 sn43_59 78000.000000
Rwneg43_60 in43_60 sn43_60 202000.000000
Rwneg43_61 in43_61 sn43_61 202000.000000
Rwneg43_62 in43_62 sn43_62 78000.000000
Rwneg43_63 in43_63 sn43_63 202000.000000
Rwneg43_64 in43_64 sn43_64 78000.000000
Rwneg43_65 in43_65 sn43_65 78000.000000
Rwneg43_66 in43_66 sn43_66 202000.000000
Rwneg43_67 in43_67 sn43_67 202000.000000
Rwneg43_68 in43_68 sn43_68 78000.000000
Rwneg43_69 in43_69 sn43_69 202000.000000
Rwneg43_70 in43_70 sn43_70 202000.000000
Rwneg43_71 in43_71 sn43_71 202000.000000
Rwneg43_72 in43_72 sn43_72 78000.000000
Rwneg43_73 in43_73 sn43_73 202000.000000
Rwneg43_74 in43_74 sn43_74 202000.000000
Rwneg43_75 in43_75 sn43_75 202000.000000
Rwneg43_76 in43_76 sn43_76 202000.000000
Rwneg43_77 in43_77 sn43_77 78000.000000
Rwneg43_78 in43_78 sn43_78 78000.000000
Rwneg43_79 in43_79 sn43_79 202000.000000
Rwneg43_80 in43_80 sn43_80 78000.000000
Rwneg43_81 in43_81 sn43_81 78000.000000
Rwneg43_82 in43_82 sn43_82 202000.000000
Rwneg43_83 in43_83 sn43_83 78000.000000
Rwneg43_84 in43_84 sn43_84 78000.000000
Rwneg44_1 in44_1 sn44_1 78000.000000
Rwneg44_2 in44_2 sn44_2 78000.000000
Rwneg44_3 in44_3 sn44_3 202000.000000
Rwneg44_4 in44_4 sn44_4 78000.000000
Rwneg44_5 in44_5 sn44_5 202000.000000
Rwneg44_6 in44_6 sn44_6 78000.000000
Rwneg44_7 in44_7 sn44_7 78000.000000
Rwneg44_8 in44_8 sn44_8 202000.000000
Rwneg44_9 in44_9 sn44_9 202000.000000
Rwneg44_10 in44_10 sn44_10 202000.000000
Rwneg44_11 in44_11 sn44_11 78000.000000
Rwneg44_12 in44_12 sn44_12 78000.000000
Rwneg44_13 in44_13 sn44_13 202000.000000
Rwneg44_14 in44_14 sn44_14 202000.000000
Rwneg44_15 in44_15 sn44_15 78000.000000
Rwneg44_16 in44_16 sn44_16 78000.000000
Rwneg44_17 in44_17 sn44_17 78000.000000
Rwneg44_18 in44_18 sn44_18 202000.000000
Rwneg44_19 in44_19 sn44_19 202000.000000
Rwneg44_20 in44_20 sn44_20 202000.000000
Rwneg44_21 in44_21 sn44_21 202000.000000
Rwneg44_22 in44_22 sn44_22 202000.000000
Rwneg44_23 in44_23 sn44_23 78000.000000
Rwneg44_24 in44_24 sn44_24 78000.000000
Rwneg44_25 in44_25 sn44_25 202000.000000
Rwneg44_26 in44_26 sn44_26 202000.000000
Rwneg44_27 in44_27 sn44_27 202000.000000
Rwneg44_28 in44_28 sn44_28 78000.000000
Rwneg44_29 in44_29 sn44_29 202000.000000
Rwneg44_30 in44_30 sn44_30 202000.000000
Rwneg44_31 in44_31 sn44_31 202000.000000
Rwneg44_32 in44_32 sn44_32 78000.000000
Rwneg44_33 in44_33 sn44_33 202000.000000
Rwneg44_34 in44_34 sn44_34 202000.000000
Rwneg44_35 in44_35 sn44_35 202000.000000
Rwneg44_36 in44_36 sn44_36 78000.000000
Rwneg44_37 in44_37 sn44_37 78000.000000
Rwneg44_38 in44_38 sn44_38 202000.000000
Rwneg44_39 in44_39 sn44_39 202000.000000
Rwneg44_40 in44_40 sn44_40 78000.000000
Rwneg44_41 in44_41 sn44_41 78000.000000
Rwneg44_42 in44_42 sn44_42 78000.000000
Rwneg44_43 in44_43 sn44_43 202000.000000
Rwneg44_44 in44_44 sn44_44 78000.000000
Rwneg44_45 in44_45 sn44_45 202000.000000
Rwneg44_46 in44_46 sn44_46 202000.000000
Rwneg44_47 in44_47 sn44_47 202000.000000
Rwneg44_48 in44_48 sn44_48 78000.000000
Rwneg44_49 in44_49 sn44_49 202000.000000
Rwneg44_50 in44_50 sn44_50 202000.000000
Rwneg44_51 in44_51 sn44_51 202000.000000
Rwneg44_52 in44_52 sn44_52 202000.000000
Rwneg44_53 in44_53 sn44_53 78000.000000
Rwneg44_54 in44_54 sn44_54 202000.000000
Rwneg44_55 in44_55 sn44_55 202000.000000
Rwneg44_56 in44_56 sn44_56 78000.000000
Rwneg44_57 in44_57 sn44_57 78000.000000
Rwneg44_58 in44_58 sn44_58 202000.000000
Rwneg44_59 in44_59 sn44_59 78000.000000
Rwneg44_60 in44_60 sn44_60 78000.000000
Rwneg44_61 in44_61 sn44_61 78000.000000
Rwneg44_62 in44_62 sn44_62 78000.000000
Rwneg44_63 in44_63 sn44_63 202000.000000
Rwneg44_64 in44_64 sn44_64 78000.000000
Rwneg44_65 in44_65 sn44_65 78000.000000
Rwneg44_66 in44_66 sn44_66 202000.000000
Rwneg44_67 in44_67 sn44_67 202000.000000
Rwneg44_68 in44_68 sn44_68 78000.000000
Rwneg44_69 in44_69 sn44_69 202000.000000
Rwneg44_70 in44_70 sn44_70 202000.000000
Rwneg44_71 in44_71 sn44_71 202000.000000
Rwneg44_72 in44_72 sn44_72 202000.000000
Rwneg44_73 in44_73 sn44_73 78000.000000
Rwneg44_74 in44_74 sn44_74 78000.000000
Rwneg44_75 in44_75 sn44_75 202000.000000
Rwneg44_76 in44_76 sn44_76 202000.000000
Rwneg44_77 in44_77 sn44_77 202000.000000
Rwneg44_78 in44_78 sn44_78 78000.000000
Rwneg44_79 in44_79 sn44_79 78000.000000
Rwneg44_80 in44_80 sn44_80 202000.000000
Rwneg44_81 in44_81 sn44_81 78000.000000
Rwneg44_82 in44_82 sn44_82 202000.000000
Rwneg44_83 in44_83 sn44_83 78000.000000
Rwneg44_84 in44_84 sn44_84 202000.000000
Rwneg45_1 in45_1 sn45_1 78000.000000
Rwneg45_2 in45_2 sn45_2 78000.000000
Rwneg45_3 in45_3 sn45_3 202000.000000
Rwneg45_4 in45_4 sn45_4 78000.000000
Rwneg45_5 in45_5 sn45_5 202000.000000
Rwneg45_6 in45_6 sn45_6 78000.000000
Rwneg45_7 in45_7 sn45_7 78000.000000
Rwneg45_8 in45_8 sn45_8 78000.000000
Rwneg45_9 in45_9 sn45_9 78000.000000
Rwneg45_10 in45_10 sn45_10 202000.000000
Rwneg45_11 in45_11 sn45_11 202000.000000
Rwneg45_12 in45_12 sn45_12 78000.000000
Rwneg45_13 in45_13 sn45_13 78000.000000
Rwneg45_14 in45_14 sn45_14 78000.000000
Rwneg45_15 in45_15 sn45_15 202000.000000
Rwneg45_16 in45_16 sn45_16 78000.000000
Rwneg45_17 in45_17 sn45_17 78000.000000
Rwneg45_18 in45_18 sn45_18 202000.000000
Rwneg45_19 in45_19 sn45_19 202000.000000
Rwneg45_20 in45_20 sn45_20 202000.000000
Rwneg45_21 in45_21 sn45_21 78000.000000
Rwneg45_22 in45_22 sn45_22 78000.000000
Rwneg45_23 in45_23 sn45_23 202000.000000
Rwneg45_24 in45_24 sn45_24 78000.000000
Rwneg45_25 in45_25 sn45_25 202000.000000
Rwneg45_26 in45_26 sn45_26 78000.000000
Rwneg45_27 in45_27 sn45_27 78000.000000
Rwneg45_28 in45_28 sn45_28 78000.000000
Rwneg45_29 in45_29 sn45_29 78000.000000
Rwneg45_30 in45_30 sn45_30 78000.000000
Rwneg45_31 in45_31 sn45_31 78000.000000
Rwneg45_32 in45_32 sn45_32 202000.000000
Rwneg45_33 in45_33 sn45_33 202000.000000
Rwneg45_34 in45_34 sn45_34 78000.000000
Rwneg45_35 in45_35 sn45_35 202000.000000
Rwneg45_36 in45_36 sn45_36 78000.000000
Rwneg45_37 in45_37 sn45_37 78000.000000
Rwneg45_38 in45_38 sn45_38 78000.000000
Rwneg45_39 in45_39 sn45_39 78000.000000
Rwneg45_40 in45_40 sn45_40 202000.000000
Rwneg45_41 in45_41 sn45_41 202000.000000
Rwneg45_42 in45_42 sn45_42 78000.000000
Rwneg45_43 in45_43 sn45_43 78000.000000
Rwneg45_44 in45_44 sn45_44 202000.000000
Rwneg45_45 in45_45 sn45_45 202000.000000
Rwneg45_46 in45_46 sn45_46 78000.000000
Rwneg45_47 in45_47 sn45_47 78000.000000
Rwneg45_48 in45_48 sn45_48 202000.000000
Rwneg45_49 in45_49 sn45_49 202000.000000
Rwneg45_50 in45_50 sn45_50 202000.000000
Rwneg45_51 in45_51 sn45_51 78000.000000
Rwneg45_52 in45_52 sn45_52 78000.000000
Rwneg45_53 in45_53 sn45_53 78000.000000
Rwneg45_54 in45_54 sn45_54 78000.000000
Rwneg45_55 in45_55 sn45_55 202000.000000
Rwneg45_56 in45_56 sn45_56 202000.000000
Rwneg45_57 in45_57 sn45_57 202000.000000
Rwneg45_58 in45_58 sn45_58 202000.000000
Rwneg45_59 in45_59 sn45_59 78000.000000
Rwneg45_60 in45_60 sn45_60 78000.000000
Rwneg45_61 in45_61 sn45_61 202000.000000
Rwneg45_62 in45_62 sn45_62 78000.000000
Rwneg45_63 in45_63 sn45_63 202000.000000
Rwneg45_64 in45_64 sn45_64 78000.000000
Rwneg45_65 in45_65 sn45_65 202000.000000
Rwneg45_66 in45_66 sn45_66 202000.000000
Rwneg45_67 in45_67 sn45_67 78000.000000
Rwneg45_68 in45_68 sn45_68 78000.000000
Rwneg45_69 in45_69 sn45_69 202000.000000
Rwneg45_70 in45_70 sn45_70 78000.000000
Rwneg45_71 in45_71 sn45_71 202000.000000
Rwneg45_72 in45_72 sn45_72 78000.000000
Rwneg45_73 in45_73 sn45_73 78000.000000
Rwneg45_74 in45_74 sn45_74 202000.000000
Rwneg45_75 in45_75 sn45_75 202000.000000
Rwneg45_76 in45_76 sn45_76 78000.000000
Rwneg45_77 in45_77 sn45_77 202000.000000
Rwneg45_78 in45_78 sn45_78 78000.000000
Rwneg45_79 in45_79 sn45_79 202000.000000
Rwneg45_80 in45_80 sn45_80 202000.000000
Rwneg45_81 in45_81 sn45_81 202000.000000
Rwneg45_82 in45_82 sn45_82 78000.000000
Rwneg45_83 in45_83 sn45_83 202000.000000
Rwneg45_84 in45_84 sn45_84 202000.000000
Rwneg46_1 in46_1 sn46_1 202000.000000
Rwneg46_2 in46_2 sn46_2 202000.000000
Rwneg46_3 in46_3 sn46_3 202000.000000
Rwneg46_4 in46_4 sn46_4 78000.000000
Rwneg46_5 in46_5 sn46_5 202000.000000
Rwneg46_6 in46_6 sn46_6 202000.000000
Rwneg46_7 in46_7 sn46_7 202000.000000
Rwneg46_8 in46_8 sn46_8 78000.000000
Rwneg46_9 in46_9 sn46_9 78000.000000
Rwneg46_10 in46_10 sn46_10 78000.000000
Rwneg46_11 in46_11 sn46_11 202000.000000
Rwneg46_12 in46_12 sn46_12 78000.000000
Rwneg46_13 in46_13 sn46_13 202000.000000
Rwneg46_14 in46_14 sn46_14 202000.000000
Rwneg46_15 in46_15 sn46_15 202000.000000
Rwneg46_16 in46_16 sn46_16 78000.000000
Rwneg46_17 in46_17 sn46_17 202000.000000
Rwneg46_18 in46_18 sn46_18 202000.000000
Rwneg46_19 in46_19 sn46_19 78000.000000
Rwneg46_20 in46_20 sn46_20 78000.000000
Rwneg46_21 in46_21 sn46_21 78000.000000
Rwneg46_22 in46_22 sn46_22 202000.000000
Rwneg46_23 in46_23 sn46_23 202000.000000
Rwneg46_24 in46_24 sn46_24 202000.000000
Rwneg46_25 in46_25 sn46_25 202000.000000
Rwneg46_26 in46_26 sn46_26 202000.000000
Rwneg46_27 in46_27 sn46_27 78000.000000
Rwneg46_28 in46_28 sn46_28 78000.000000
Rwneg46_29 in46_29 sn46_29 78000.000000
Rwneg46_30 in46_30 sn46_30 78000.000000
Rwneg46_31 in46_31 sn46_31 202000.000000
Rwneg46_32 in46_32 sn46_32 202000.000000
Rwneg46_33 in46_33 sn46_33 202000.000000
Rwneg46_34 in46_34 sn46_34 78000.000000
Rwneg46_35 in46_35 sn46_35 202000.000000
Rwneg46_36 in46_36 sn46_36 202000.000000
Rwneg46_37 in46_37 sn46_37 78000.000000
Rwneg46_38 in46_38 sn46_38 202000.000000
Rwneg46_39 in46_39 sn46_39 202000.000000
Rwneg46_40 in46_40 sn46_40 78000.000000
Rwneg46_41 in46_41 sn46_41 202000.000000
Rwneg46_42 in46_42 sn46_42 202000.000000
Rwneg46_43 in46_43 sn46_43 78000.000000
Rwneg46_44 in46_44 sn46_44 78000.000000
Rwneg46_45 in46_45 sn46_45 78000.000000
Rwneg46_46 in46_46 sn46_46 202000.000000
Rwneg46_47 in46_47 sn46_47 202000.000000
Rwneg46_48 in46_48 sn46_48 78000.000000
Rwneg46_49 in46_49 sn46_49 78000.000000
Rwneg46_50 in46_50 sn46_50 78000.000000
Rwneg46_51 in46_51 sn46_51 202000.000000
Rwneg46_52 in46_52 sn46_52 78000.000000
Rwneg46_53 in46_53 sn46_53 78000.000000
Rwneg46_54 in46_54 sn46_54 78000.000000
Rwneg46_55 in46_55 sn46_55 78000.000000
Rwneg46_56 in46_56 sn46_56 202000.000000
Rwneg46_57 in46_57 sn46_57 202000.000000
Rwneg46_58 in46_58 sn46_58 202000.000000
Rwneg46_59 in46_59 sn46_59 202000.000000
Rwneg46_60 in46_60 sn46_60 78000.000000
Rwneg46_61 in46_61 sn46_61 202000.000000
Rwneg46_62 in46_62 sn46_62 202000.000000
Rwneg46_63 in46_63 sn46_63 78000.000000
Rwneg46_64 in46_64 sn46_64 78000.000000
Rwneg46_65 in46_65 sn46_65 202000.000000
Rwneg46_66 in46_66 sn46_66 78000.000000
Rwneg46_67 in46_67 sn46_67 202000.000000
Rwneg46_68 in46_68 sn46_68 78000.000000
Rwneg46_69 in46_69 sn46_69 78000.000000
Rwneg46_70 in46_70 sn46_70 202000.000000
Rwneg46_71 in46_71 sn46_71 78000.000000
Rwneg46_72 in46_72 sn46_72 202000.000000
Rwneg46_73 in46_73 sn46_73 78000.000000
Rwneg46_74 in46_74 sn46_74 202000.000000
Rwneg46_75 in46_75 sn46_75 202000.000000
Rwneg46_76 in46_76 sn46_76 202000.000000
Rwneg46_77 in46_77 sn46_77 202000.000000
Rwneg46_78 in46_78 sn46_78 78000.000000
Rwneg46_79 in46_79 sn46_79 202000.000000
Rwneg46_80 in46_80 sn46_80 202000.000000
Rwneg46_81 in46_81 sn46_81 202000.000000
Rwneg46_82 in46_82 sn46_82 78000.000000
Rwneg46_83 in46_83 sn46_83 202000.000000
Rwneg46_84 in46_84 sn46_84 202000.000000
Rwneg47_1 in47_1 sn47_1 202000.000000
Rwneg47_2 in47_2 sn47_2 202000.000000
Rwneg47_3 in47_3 sn47_3 78000.000000
Rwneg47_4 in47_4 sn47_4 78000.000000
Rwneg47_5 in47_5 sn47_5 78000.000000
Rwneg47_6 in47_6 sn47_6 78000.000000
Rwneg47_7 in47_7 sn47_7 202000.000000
Rwneg47_8 in47_8 sn47_8 202000.000000
Rwneg47_9 in47_9 sn47_9 202000.000000
Rwneg47_10 in47_10 sn47_10 202000.000000
Rwneg47_11 in47_11 sn47_11 202000.000000
Rwneg47_12 in47_12 sn47_12 202000.000000
Rwneg47_13 in47_13 sn47_13 78000.000000
Rwneg47_14 in47_14 sn47_14 202000.000000
Rwneg47_15 in47_15 sn47_15 202000.000000
Rwneg47_16 in47_16 sn47_16 202000.000000
Rwneg47_17 in47_17 sn47_17 78000.000000
Rwneg47_18 in47_18 sn47_18 202000.000000
Rwneg47_19 in47_19 sn47_19 202000.000000
Rwneg47_20 in47_20 sn47_20 202000.000000
Rwneg47_21 in47_21 sn47_21 202000.000000
Rwneg47_22 in47_22 sn47_22 78000.000000
Rwneg47_23 in47_23 sn47_23 202000.000000
Rwneg47_24 in47_24 sn47_24 78000.000000
Rwneg47_25 in47_25 sn47_25 78000.000000
Rwneg47_26 in47_26 sn47_26 202000.000000
Rwneg47_27 in47_27 sn47_27 78000.000000
Rwneg47_28 in47_28 sn47_28 202000.000000
Rwneg47_29 in47_29 sn47_29 78000.000000
Rwneg47_30 in47_30 sn47_30 78000.000000
Rwneg47_31 in47_31 sn47_31 78000.000000
Rwneg47_32 in47_32 sn47_32 202000.000000
Rwneg47_33 in47_33 sn47_33 202000.000000
Rwneg47_34 in47_34 sn47_34 202000.000000
Rwneg47_35 in47_35 sn47_35 78000.000000
Rwneg47_36 in47_36 sn47_36 202000.000000
Rwneg47_37 in47_37 sn47_37 202000.000000
Rwneg47_38 in47_38 sn47_38 202000.000000
Rwneg47_39 in47_39 sn47_39 78000.000000
Rwneg47_40 in47_40 sn47_40 202000.000000
Rwneg47_41 in47_41 sn47_41 78000.000000
Rwneg47_42 in47_42 sn47_42 202000.000000
Rwneg47_43 in47_43 sn47_43 202000.000000
Rwneg47_44 in47_44 sn47_44 202000.000000
Rwneg47_45 in47_45 sn47_45 202000.000000
Rwneg47_46 in47_46 sn47_46 78000.000000
Rwneg47_47 in47_47 sn47_47 78000.000000
Rwneg47_48 in47_48 sn47_48 202000.000000
Rwneg47_49 in47_49 sn47_49 202000.000000
Rwneg47_50 in47_50 sn47_50 202000.000000
Rwneg47_51 in47_51 sn47_51 202000.000000
Rwneg47_52 in47_52 sn47_52 202000.000000
Rwneg47_53 in47_53 sn47_53 78000.000000
Rwneg47_54 in47_54 sn47_54 78000.000000
Rwneg47_55 in47_55 sn47_55 78000.000000
Rwneg47_56 in47_56 sn47_56 202000.000000
Rwneg47_57 in47_57 sn47_57 78000.000000
Rwneg47_58 in47_58 sn47_58 202000.000000
Rwneg47_59 in47_59 sn47_59 202000.000000
Rwneg47_60 in47_60 sn47_60 202000.000000
Rwneg47_61 in47_61 sn47_61 202000.000000
Rwneg47_62 in47_62 sn47_62 78000.000000
Rwneg47_63 in47_63 sn47_63 202000.000000
Rwneg47_64 in47_64 sn47_64 78000.000000
Rwneg47_65 in47_65 sn47_65 78000.000000
Rwneg47_66 in47_66 sn47_66 202000.000000
Rwneg47_67 in47_67 sn47_67 202000.000000
Rwneg47_68 in47_68 sn47_68 78000.000000
Rwneg47_69 in47_69 sn47_69 202000.000000
Rwneg47_70 in47_70 sn47_70 78000.000000
Rwneg47_71 in47_71 sn47_71 202000.000000
Rwneg47_72 in47_72 sn47_72 202000.000000
Rwneg47_73 in47_73 sn47_73 202000.000000
Rwneg47_74 in47_74 sn47_74 78000.000000
Rwneg47_75 in47_75 sn47_75 78000.000000
Rwneg47_76 in47_76 sn47_76 202000.000000
Rwneg47_77 in47_77 sn47_77 202000.000000
Rwneg47_78 in47_78 sn47_78 202000.000000
Rwneg47_79 in47_79 sn47_79 202000.000000
Rwneg47_80 in47_80 sn47_80 78000.000000
Rwneg47_81 in47_81 sn47_81 78000.000000
Rwneg47_82 in47_82 sn47_82 202000.000000
Rwneg47_83 in47_83 sn47_83 202000.000000
Rwneg47_84 in47_84 sn47_84 202000.000000
Rwneg48_1 in48_1 sn48_1 202000.000000
Rwneg48_2 in48_2 sn48_2 78000.000000
Rwneg48_3 in48_3 sn48_3 202000.000000
Rwneg48_4 in48_4 sn48_4 202000.000000
Rwneg48_5 in48_5 sn48_5 78000.000000
Rwneg48_6 in48_6 sn48_6 78000.000000
Rwneg48_7 in48_7 sn48_7 78000.000000
Rwneg48_8 in48_8 sn48_8 78000.000000
Rwneg48_9 in48_9 sn48_9 202000.000000
Rwneg48_10 in48_10 sn48_10 202000.000000
Rwneg48_11 in48_11 sn48_11 202000.000000
Rwneg48_12 in48_12 sn48_12 202000.000000
Rwneg48_13 in48_13 sn48_13 202000.000000
Rwneg48_14 in48_14 sn48_14 78000.000000
Rwneg48_15 in48_15 sn48_15 78000.000000
Rwneg48_16 in48_16 sn48_16 78000.000000
Rwneg48_17 in48_17 sn48_17 202000.000000
Rwneg48_18 in48_18 sn48_18 78000.000000
Rwneg48_19 in48_19 sn48_19 202000.000000
Rwneg48_20 in48_20 sn48_20 78000.000000
Rwneg48_21 in48_21 sn48_21 78000.000000
Rwneg48_22 in48_22 sn48_22 202000.000000
Rwneg48_23 in48_23 sn48_23 202000.000000
Rwneg48_24 in48_24 sn48_24 78000.000000
Rwneg48_25 in48_25 sn48_25 202000.000000
Rwneg48_26 in48_26 sn48_26 202000.000000
Rwneg48_27 in48_27 sn48_27 202000.000000
Rwneg48_28 in48_28 sn48_28 202000.000000
Rwneg48_29 in48_29 sn48_29 78000.000000
Rwneg48_30 in48_30 sn48_30 202000.000000
Rwneg48_31 in48_31 sn48_31 202000.000000
Rwneg48_32 in48_32 sn48_32 202000.000000
Rwneg48_33 in48_33 sn48_33 202000.000000
Rwneg48_34 in48_34 sn48_34 202000.000000
Rwneg48_35 in48_35 sn48_35 202000.000000
Rwneg48_36 in48_36 sn48_36 78000.000000
Rwneg48_37 in48_37 sn48_37 202000.000000
Rwneg48_38 in48_38 sn48_38 78000.000000
Rwneg48_39 in48_39 sn48_39 202000.000000
Rwneg48_40 in48_40 sn48_40 202000.000000
Rwneg48_41 in48_41 sn48_41 202000.000000
Rwneg48_42 in48_42 sn48_42 78000.000000
Rwneg48_43 in48_43 sn48_43 78000.000000
Rwneg48_44 in48_44 sn48_44 78000.000000
Rwneg48_45 in48_45 sn48_45 78000.000000
Rwneg48_46 in48_46 sn48_46 202000.000000
Rwneg48_47 in48_47 sn48_47 78000.000000
Rwneg48_48 in48_48 sn48_48 202000.000000
Rwneg48_49 in48_49 sn48_49 78000.000000
Rwneg48_50 in48_50 sn48_50 78000.000000
Rwneg48_51 in48_51 sn48_51 202000.000000
Rwneg48_52 in48_52 sn48_52 78000.000000
Rwneg48_53 in48_53 sn48_53 78000.000000
Rwneg48_54 in48_54 sn48_54 78000.000000
Rwneg48_55 in48_55 sn48_55 202000.000000
Rwneg48_56 in48_56 sn48_56 202000.000000
Rwneg48_57 in48_57 sn48_57 202000.000000
Rwneg48_58 in48_58 sn48_58 202000.000000
Rwneg48_59 in48_59 sn48_59 202000.000000
Rwneg48_60 in48_60 sn48_60 78000.000000
Rwneg48_61 in48_61 sn48_61 202000.000000
Rwneg48_62 in48_62 sn48_62 202000.000000
Rwneg48_63 in48_63 sn48_63 78000.000000
Rwneg48_64 in48_64 sn48_64 78000.000000
Rwneg48_65 in48_65 sn48_65 78000.000000
Rwneg48_66 in48_66 sn48_66 202000.000000
Rwneg48_67 in48_67 sn48_67 202000.000000
Rwneg48_68 in48_68 sn48_68 78000.000000
Rwneg48_69 in48_69 sn48_69 202000.000000
Rwneg48_70 in48_70 sn48_70 202000.000000
Rwneg48_71 in48_71 sn48_71 202000.000000
Rwneg48_72 in48_72 sn48_72 202000.000000
Rwneg48_73 in48_73 sn48_73 202000.000000
Rwneg48_74 in48_74 sn48_74 202000.000000
Rwneg48_75 in48_75 sn48_75 202000.000000
Rwneg48_76 in48_76 sn48_76 78000.000000
Rwneg48_77 in48_77 sn48_77 202000.000000
Rwneg48_78 in48_78 sn48_78 78000.000000
Rwneg48_79 in48_79 sn48_79 202000.000000
Rwneg48_80 in48_80 sn48_80 202000.000000
Rwneg48_81 in48_81 sn48_81 78000.000000
Rwneg48_82 in48_82 sn48_82 78000.000000
Rwneg48_83 in48_83 sn48_83 78000.000000
Rwneg48_84 in48_84 sn48_84 78000.000000
Rwneg49_1 in49_1 sn49_1 202000.000000
Rwneg49_2 in49_2 sn49_2 78000.000000
Rwneg49_3 in49_3 sn49_3 202000.000000
Rwneg49_4 in49_4 sn49_4 78000.000000
Rwneg49_5 in49_5 sn49_5 202000.000000
Rwneg49_6 in49_6 sn49_6 78000.000000
Rwneg49_7 in49_7 sn49_7 78000.000000
Rwneg49_8 in49_8 sn49_8 202000.000000
Rwneg49_9 in49_9 sn49_9 202000.000000
Rwneg49_10 in49_10 sn49_10 202000.000000
Rwneg49_11 in49_11 sn49_11 78000.000000
Rwneg49_12 in49_12 sn49_12 202000.000000
Rwneg49_13 in49_13 sn49_13 202000.000000
Rwneg49_14 in49_14 sn49_14 202000.000000
Rwneg49_15 in49_15 sn49_15 202000.000000
Rwneg49_16 in49_16 sn49_16 202000.000000
Rwneg49_17 in49_17 sn49_17 78000.000000
Rwneg49_18 in49_18 sn49_18 202000.000000
Rwneg49_19 in49_19 sn49_19 202000.000000
Rwneg49_20 in49_20 sn49_20 202000.000000
Rwneg49_21 in49_21 sn49_21 202000.000000
Rwneg49_22 in49_22 sn49_22 202000.000000
Rwneg49_23 in49_23 sn49_23 202000.000000
Rwneg49_24 in49_24 sn49_24 78000.000000
Rwneg49_25 in49_25 sn49_25 78000.000000
Rwneg49_26 in49_26 sn49_26 78000.000000
Rwneg49_27 in49_27 sn49_27 202000.000000
Rwneg49_28 in49_28 sn49_28 202000.000000
Rwneg49_29 in49_29 sn49_29 202000.000000
Rwneg49_30 in49_30 sn49_30 78000.000000
Rwneg49_31 in49_31 sn49_31 202000.000000
Rwneg49_32 in49_32 sn49_32 78000.000000
Rwneg49_33 in49_33 sn49_33 202000.000000
Rwneg49_34 in49_34 sn49_34 78000.000000
Rwneg49_35 in49_35 sn49_35 202000.000000
Rwneg49_36 in49_36 sn49_36 202000.000000
Rwneg49_37 in49_37 sn49_37 78000.000000
Rwneg49_38 in49_38 sn49_38 202000.000000
Rwneg49_39 in49_39 sn49_39 202000.000000
Rwneg49_40 in49_40 sn49_40 202000.000000
Rwneg49_41 in49_41 sn49_41 202000.000000
Rwneg49_42 in49_42 sn49_42 78000.000000
Rwneg49_43 in49_43 sn49_43 202000.000000
Rwneg49_44 in49_44 sn49_44 78000.000000
Rwneg49_45 in49_45 sn49_45 202000.000000
Rwneg49_46 in49_46 sn49_46 78000.000000
Rwneg49_47 in49_47 sn49_47 78000.000000
Rwneg49_48 in49_48 sn49_48 78000.000000
Rwneg49_49 in49_49 sn49_49 202000.000000
Rwneg49_50 in49_50 sn49_50 78000.000000
Rwneg49_51 in49_51 sn49_51 78000.000000
Rwneg49_52 in49_52 sn49_52 202000.000000
Rwneg49_53 in49_53 sn49_53 78000.000000
Rwneg49_54 in49_54 sn49_54 202000.000000
Rwneg49_55 in49_55 sn49_55 78000.000000
Rwneg49_56 in49_56 sn49_56 78000.000000
Rwneg49_57 in49_57 sn49_57 202000.000000
Rwneg49_58 in49_58 sn49_58 202000.000000
Rwneg49_59 in49_59 sn49_59 202000.000000
Rwneg49_60 in49_60 sn49_60 78000.000000
Rwneg49_61 in49_61 sn49_61 202000.000000
Rwneg49_62 in49_62 sn49_62 78000.000000
Rwneg49_63 in49_63 sn49_63 78000.000000
Rwneg49_64 in49_64 sn49_64 78000.000000
Rwneg49_65 in49_65 sn49_65 78000.000000
Rwneg49_66 in49_66 sn49_66 202000.000000
Rwneg49_67 in49_67 sn49_67 202000.000000
Rwneg49_68 in49_68 sn49_68 78000.000000
Rwneg49_69 in49_69 sn49_69 78000.000000
Rwneg49_70 in49_70 sn49_70 202000.000000
Rwneg49_71 in49_71 sn49_71 78000.000000
Rwneg49_72 in49_72 sn49_72 202000.000000
Rwneg49_73 in49_73 sn49_73 202000.000000
Rwneg49_74 in49_74 sn49_74 202000.000000
Rwneg49_75 in49_75 sn49_75 202000.000000
Rwneg49_76 in49_76 sn49_76 202000.000000
Rwneg49_77 in49_77 sn49_77 78000.000000
Rwneg49_78 in49_78 sn49_78 78000.000000
Rwneg49_79 in49_79 sn49_79 78000.000000
Rwneg49_80 in49_80 sn49_80 78000.000000
Rwneg49_81 in49_81 sn49_81 78000.000000
Rwneg49_82 in49_82 sn49_82 202000.000000
Rwneg49_83 in49_83 sn49_83 202000.000000
Rwneg49_84 in49_84 sn49_84 78000.000000
Rwneg50_1 in50_1 sn50_1 202000.000000
Rwneg50_2 in50_2 sn50_2 202000.000000
Rwneg50_3 in50_3 sn50_3 202000.000000
Rwneg50_4 in50_4 sn50_4 78000.000000
Rwneg50_5 in50_5 sn50_5 202000.000000
Rwneg50_6 in50_6 sn50_6 202000.000000
Rwneg50_7 in50_7 sn50_7 78000.000000
Rwneg50_8 in50_8 sn50_8 202000.000000
Rwneg50_9 in50_9 sn50_9 202000.000000
Rwneg50_10 in50_10 sn50_10 202000.000000
Rwneg50_11 in50_11 sn50_11 202000.000000
Rwneg50_12 in50_12 sn50_12 78000.000000
Rwneg50_13 in50_13 sn50_13 202000.000000
Rwneg50_14 in50_14 sn50_14 202000.000000
Rwneg50_15 in50_15 sn50_15 202000.000000
Rwneg50_16 in50_16 sn50_16 78000.000000
Rwneg50_17 in50_17 sn50_17 202000.000000
Rwneg50_18 in50_18 sn50_18 78000.000000
Rwneg50_19 in50_19 sn50_19 78000.000000
Rwneg50_20 in50_20 sn50_20 202000.000000
Rwneg50_21 in50_21 sn50_21 202000.000000
Rwneg50_22 in50_22 sn50_22 202000.000000
Rwneg50_23 in50_23 sn50_23 78000.000000
Rwneg50_24 in50_24 sn50_24 202000.000000
Rwneg50_25 in50_25 sn50_25 202000.000000
Rwneg50_26 in50_26 sn50_26 202000.000000
Rwneg50_27 in50_27 sn50_27 202000.000000
Rwneg50_28 in50_28 sn50_28 78000.000000
Rwneg50_29 in50_29 sn50_29 78000.000000
Rwneg50_30 in50_30 sn50_30 202000.000000
Rwneg50_31 in50_31 sn50_31 202000.000000
Rwneg50_32 in50_32 sn50_32 202000.000000
Rwneg50_33 in50_33 sn50_33 202000.000000
Rwneg50_34 in50_34 sn50_34 202000.000000
Rwneg50_35 in50_35 sn50_35 202000.000000
Rwneg50_36 in50_36 sn50_36 202000.000000
Rwneg50_37 in50_37 sn50_37 78000.000000
Rwneg50_38 in50_38 sn50_38 78000.000000
Rwneg50_39 in50_39 sn50_39 78000.000000
Rwneg50_40 in50_40 sn50_40 78000.000000
Rwneg50_41 in50_41 sn50_41 202000.000000
Rwneg50_42 in50_42 sn50_42 78000.000000
Rwneg50_43 in50_43 sn50_43 78000.000000
Rwneg50_44 in50_44 sn50_44 78000.000000
Rwneg50_45 in50_45 sn50_45 202000.000000
Rwneg50_46 in50_46 sn50_46 202000.000000
Rwneg50_47 in50_47 sn50_47 78000.000000
Rwneg50_48 in50_48 sn50_48 78000.000000
Rwneg50_49 in50_49 sn50_49 202000.000000
Rwneg50_50 in50_50 sn50_50 202000.000000
Rwneg50_51 in50_51 sn50_51 78000.000000
Rwneg50_52 in50_52 sn50_52 202000.000000
Rwneg50_53 in50_53 sn50_53 202000.000000
Rwneg50_54 in50_54 sn50_54 78000.000000
Rwneg50_55 in50_55 sn50_55 202000.000000
Rwneg50_56 in50_56 sn50_56 78000.000000
Rwneg50_57 in50_57 sn50_57 202000.000000
Rwneg50_58 in50_58 sn50_58 202000.000000
Rwneg50_59 in50_59 sn50_59 202000.000000
Rwneg50_60 in50_60 sn50_60 78000.000000
Rwneg50_61 in50_61 sn50_61 202000.000000
Rwneg50_62 in50_62 sn50_62 78000.000000
Rwneg50_63 in50_63 sn50_63 202000.000000
Rwneg50_64 in50_64 sn50_64 202000.000000
Rwneg50_65 in50_65 sn50_65 78000.000000
Rwneg50_66 in50_66 sn50_66 78000.000000
Rwneg50_67 in50_67 sn50_67 202000.000000
Rwneg50_68 in50_68 sn50_68 78000.000000
Rwneg50_69 in50_69 sn50_69 78000.000000
Rwneg50_70 in50_70 sn50_70 202000.000000
Rwneg50_71 in50_71 sn50_71 78000.000000
Rwneg50_72 in50_72 sn50_72 202000.000000
Rwneg50_73 in50_73 sn50_73 202000.000000
Rwneg50_74 in50_74 sn50_74 202000.000000
Rwneg50_75 in50_75 sn50_75 202000.000000
Rwneg50_76 in50_76 sn50_76 202000.000000
Rwneg50_77 in50_77 sn50_77 78000.000000
Rwneg50_78 in50_78 sn50_78 202000.000000
Rwneg50_79 in50_79 sn50_79 78000.000000
Rwneg50_80 in50_80 sn50_80 202000.000000
Rwneg50_81 in50_81 sn50_81 78000.000000
Rwneg50_82 in50_82 sn50_82 202000.000000
Rwneg50_83 in50_83 sn50_83 202000.000000
Rwneg50_84 in50_84 sn50_84 202000.000000
Rwneg51_1 in51_1 sn51_1 202000.000000
Rwneg51_2 in51_2 sn51_2 202000.000000
Rwneg51_3 in51_3 sn51_3 78000.000000
Rwneg51_4 in51_4 sn51_4 202000.000000
Rwneg51_5 in51_5 sn51_5 78000.000000
Rwneg51_6 in51_6 sn51_6 202000.000000
Rwneg51_7 in51_7 sn51_7 78000.000000
Rwneg51_8 in51_8 sn51_8 78000.000000
Rwneg51_9 in51_9 sn51_9 78000.000000
Rwneg51_10 in51_10 sn51_10 202000.000000
Rwneg51_11 in51_11 sn51_11 78000.000000
Rwneg51_12 in51_12 sn51_12 202000.000000
Rwneg51_13 in51_13 sn51_13 78000.000000
Rwneg51_14 in51_14 sn51_14 202000.000000
Rwneg51_15 in51_15 sn51_15 202000.000000
Rwneg51_16 in51_16 sn51_16 202000.000000
Rwneg51_17 in51_17 sn51_17 202000.000000
Rwneg51_18 in51_18 sn51_18 78000.000000
Rwneg51_19 in51_19 sn51_19 202000.000000
Rwneg51_20 in51_20 sn51_20 78000.000000
Rwneg51_21 in51_21 sn51_21 202000.000000
Rwneg51_22 in51_22 sn51_22 202000.000000
Rwneg51_23 in51_23 sn51_23 78000.000000
Rwneg51_24 in51_24 sn51_24 202000.000000
Rwneg51_25 in51_25 sn51_25 78000.000000
Rwneg51_26 in51_26 sn51_26 202000.000000
Rwneg51_27 in51_27 sn51_27 78000.000000
Rwneg51_28 in51_28 sn51_28 202000.000000
Rwneg51_29 in51_29 sn51_29 78000.000000
Rwneg51_30 in51_30 sn51_30 202000.000000
Rwneg51_31 in51_31 sn51_31 202000.000000
Rwneg51_32 in51_32 sn51_32 78000.000000
Rwneg51_33 in51_33 sn51_33 202000.000000
Rwneg51_34 in51_34 sn51_34 78000.000000
Rwneg51_35 in51_35 sn51_35 78000.000000
Rwneg51_36 in51_36 sn51_36 78000.000000
Rwneg51_37 in51_37 sn51_37 78000.000000
Rwneg51_38 in51_38 sn51_38 202000.000000
Rwneg51_39 in51_39 sn51_39 202000.000000
Rwneg51_40 in51_40 sn51_40 202000.000000
Rwneg51_41 in51_41 sn51_41 78000.000000
Rwneg51_42 in51_42 sn51_42 78000.000000
Rwneg51_43 in51_43 sn51_43 78000.000000
Rwneg51_44 in51_44 sn51_44 202000.000000
Rwneg51_45 in51_45 sn51_45 202000.000000
Rwneg51_46 in51_46 sn51_46 78000.000000
Rwneg51_47 in51_47 sn51_47 202000.000000
Rwneg51_48 in51_48 sn51_48 78000.000000
Rwneg51_49 in51_49 sn51_49 78000.000000
Rwneg51_50 in51_50 sn51_50 202000.000000
Rwneg51_51 in51_51 sn51_51 202000.000000
Rwneg51_52 in51_52 sn51_52 202000.000000
Rwneg51_53 in51_53 sn51_53 202000.000000
Rwneg51_54 in51_54 sn51_54 202000.000000
Rwneg51_55 in51_55 sn51_55 78000.000000
Rwneg51_56 in51_56 sn51_56 78000.000000
Rwneg51_57 in51_57 sn51_57 202000.000000
Rwneg51_58 in51_58 sn51_58 78000.000000
Rwneg51_59 in51_59 sn51_59 78000.000000
Rwneg51_60 in51_60 sn51_60 78000.000000
Rwneg51_61 in51_61 sn51_61 202000.000000
Rwneg51_62 in51_62 sn51_62 78000.000000
Rwneg51_63 in51_63 sn51_63 202000.000000
Rwneg51_64 in51_64 sn51_64 78000.000000
Rwneg51_65 in51_65 sn51_65 78000.000000
Rwneg51_66 in51_66 sn51_66 78000.000000
Rwneg51_67 in51_67 sn51_67 202000.000000
Rwneg51_68 in51_68 sn51_68 202000.000000
Rwneg51_69 in51_69 sn51_69 78000.000000
Rwneg51_70 in51_70 sn51_70 202000.000000
Rwneg51_71 in51_71 sn51_71 78000.000000
Rwneg51_72 in51_72 sn51_72 202000.000000
Rwneg51_73 in51_73 sn51_73 202000.000000
Rwneg51_74 in51_74 sn51_74 202000.000000
Rwneg51_75 in51_75 sn51_75 78000.000000
Rwneg51_76 in51_76 sn51_76 78000.000000
Rwneg51_77 in51_77 sn51_77 202000.000000
Rwneg51_78 in51_78 sn51_78 202000.000000
Rwneg51_79 in51_79 sn51_79 78000.000000
Rwneg51_80 in51_80 sn51_80 78000.000000
Rwneg51_81 in51_81 sn51_81 78000.000000
Rwneg51_82 in51_82 sn51_82 202000.000000
Rwneg51_83 in51_83 sn51_83 202000.000000
Rwneg51_84 in51_84 sn51_84 202000.000000
Rwneg52_1 in52_1 sn52_1 78000.000000
Rwneg52_2 in52_2 sn52_2 78000.000000
Rwneg52_3 in52_3 sn52_3 202000.000000
Rwneg52_4 in52_4 sn52_4 202000.000000
Rwneg52_5 in52_5 sn52_5 78000.000000
Rwneg52_6 in52_6 sn52_6 78000.000000
Rwneg52_7 in52_7 sn52_7 78000.000000
Rwneg52_8 in52_8 sn52_8 202000.000000
Rwneg52_9 in52_9 sn52_9 202000.000000
Rwneg52_10 in52_10 sn52_10 78000.000000
Rwneg52_11 in52_11 sn52_11 202000.000000
Rwneg52_12 in52_12 sn52_12 202000.000000
Rwneg52_13 in52_13 sn52_13 202000.000000
Rwneg52_14 in52_14 sn52_14 78000.000000
Rwneg52_15 in52_15 sn52_15 202000.000000
Rwneg52_16 in52_16 sn52_16 202000.000000
Rwneg52_17 in52_17 sn52_17 202000.000000
Rwneg52_18 in52_18 sn52_18 78000.000000
Rwneg52_19 in52_19 sn52_19 202000.000000
Rwneg52_20 in52_20 sn52_20 202000.000000
Rwneg52_21 in52_21 sn52_21 78000.000000
Rwneg52_22 in52_22 sn52_22 202000.000000
Rwneg52_23 in52_23 sn52_23 202000.000000
Rwneg52_24 in52_24 sn52_24 78000.000000
Rwneg52_25 in52_25 sn52_25 202000.000000
Rwneg52_26 in52_26 sn52_26 202000.000000
Rwneg52_27 in52_27 sn52_27 78000.000000
Rwneg52_28 in52_28 sn52_28 202000.000000
Rwneg52_29 in52_29 sn52_29 78000.000000
Rwneg52_30 in52_30 sn52_30 202000.000000
Rwneg52_31 in52_31 sn52_31 202000.000000
Rwneg52_32 in52_32 sn52_32 78000.000000
Rwneg52_33 in52_33 sn52_33 202000.000000
Rwneg52_34 in52_34 sn52_34 78000.000000
Rwneg52_35 in52_35 sn52_35 202000.000000
Rwneg52_36 in52_36 sn52_36 78000.000000
Rwneg52_37 in52_37 sn52_37 78000.000000
Rwneg52_38 in52_38 sn52_38 202000.000000
Rwneg52_39 in52_39 sn52_39 202000.000000
Rwneg52_40 in52_40 sn52_40 202000.000000
Rwneg52_41 in52_41 sn52_41 202000.000000
Rwneg52_42 in52_42 sn52_42 78000.000000
Rwneg52_43 in52_43 sn52_43 202000.000000
Rwneg52_44 in52_44 sn52_44 78000.000000
Rwneg52_45 in52_45 sn52_45 202000.000000
Rwneg52_46 in52_46 sn52_46 78000.000000
Rwneg52_47 in52_47 sn52_47 78000.000000
Rwneg52_48 in52_48 sn52_48 78000.000000
Rwneg52_49 in52_49 sn52_49 202000.000000
Rwneg52_50 in52_50 sn52_50 78000.000000
Rwneg52_51 in52_51 sn52_51 202000.000000
Rwneg52_52 in52_52 sn52_52 78000.000000
Rwneg52_53 in52_53 sn52_53 202000.000000
Rwneg52_54 in52_54 sn52_54 78000.000000
Rwneg52_55 in52_55 sn52_55 78000.000000
Rwneg52_56 in52_56 sn52_56 202000.000000
Rwneg52_57 in52_57 sn52_57 202000.000000
Rwneg52_58 in52_58 sn52_58 202000.000000
Rwneg52_59 in52_59 sn52_59 202000.000000
Rwneg52_60 in52_60 sn52_60 78000.000000
Rwneg52_61 in52_61 sn52_61 202000.000000
Rwneg52_62 in52_62 sn52_62 78000.000000
Rwneg52_63 in52_63 sn52_63 202000.000000
Rwneg52_64 in52_64 sn52_64 202000.000000
Rwneg52_65 in52_65 sn52_65 78000.000000
Rwneg52_66 in52_66 sn52_66 78000.000000
Rwneg52_67 in52_67 sn52_67 78000.000000
Rwneg52_68 in52_68 sn52_68 78000.000000
Rwneg52_69 in52_69 sn52_69 78000.000000
Rwneg52_70 in52_70 sn52_70 202000.000000
Rwneg52_71 in52_71 sn52_71 78000.000000
Rwneg52_72 in52_72 sn52_72 202000.000000
Rwneg52_73 in52_73 sn52_73 78000.000000
Rwneg52_74 in52_74 sn52_74 202000.000000
Rwneg52_75 in52_75 sn52_75 202000.000000
Rwneg52_76 in52_76 sn52_76 202000.000000
Rwneg52_77 in52_77 sn52_77 78000.000000
Rwneg52_78 in52_78 sn52_78 202000.000000
Rwneg52_79 in52_79 sn52_79 78000.000000
Rwneg52_80 in52_80 sn52_80 202000.000000
Rwneg52_81 in52_81 sn52_81 78000.000000
Rwneg52_82 in52_82 sn52_82 78000.000000
Rwneg52_83 in52_83 sn52_83 202000.000000
Rwneg52_84 in52_84 sn52_84 202000.000000
Rwneg53_1 in53_1 sn53_1 202000.000000
Rwneg53_2 in53_2 sn53_2 78000.000000
Rwneg53_3 in53_3 sn53_3 202000.000000
Rwneg53_4 in53_4 sn53_4 78000.000000
Rwneg53_5 in53_5 sn53_5 78000.000000
Rwneg53_6 in53_6 sn53_6 202000.000000
Rwneg53_7 in53_7 sn53_7 202000.000000
Rwneg53_8 in53_8 sn53_8 78000.000000
Rwneg53_9 in53_9 sn53_9 78000.000000
Rwneg53_10 in53_10 sn53_10 202000.000000
Rwneg53_11 in53_11 sn53_11 78000.000000
Rwneg53_12 in53_12 sn53_12 78000.000000
Rwneg53_13 in53_13 sn53_13 202000.000000
Rwneg53_14 in53_14 sn53_14 78000.000000
Rwneg53_15 in53_15 sn53_15 202000.000000
Rwneg53_16 in53_16 sn53_16 78000.000000
Rwneg53_17 in53_17 sn53_17 202000.000000
Rwneg53_18 in53_18 sn53_18 202000.000000
Rwneg53_19 in53_19 sn53_19 202000.000000
Rwneg53_20 in53_20 sn53_20 202000.000000
Rwneg53_21 in53_21 sn53_21 202000.000000
Rwneg53_22 in53_22 sn53_22 78000.000000
Rwneg53_23 in53_23 sn53_23 202000.000000
Rwneg53_24 in53_24 sn53_24 202000.000000
Rwneg53_25 in53_25 sn53_25 78000.000000
Rwneg53_26 in53_26 sn53_26 202000.000000
Rwneg53_27 in53_27 sn53_27 78000.000000
Rwneg53_28 in53_28 sn53_28 202000.000000
Rwneg53_29 in53_29 sn53_29 202000.000000
Rwneg53_30 in53_30 sn53_30 78000.000000
Rwneg53_31 in53_31 sn53_31 78000.000000
Rwneg53_32 in53_32 sn53_32 202000.000000
Rwneg53_33 in53_33 sn53_33 202000.000000
Rwneg53_34 in53_34 sn53_34 78000.000000
Rwneg53_35 in53_35 sn53_35 78000.000000
Rwneg53_36 in53_36 sn53_36 78000.000000
Rwneg53_37 in53_37 sn53_37 202000.000000
Rwneg53_38 in53_38 sn53_38 202000.000000
Rwneg53_39 in53_39 sn53_39 202000.000000
Rwneg53_40 in53_40 sn53_40 202000.000000
Rwneg53_41 in53_41 sn53_41 78000.000000
Rwneg53_42 in53_42 sn53_42 202000.000000
Rwneg53_43 in53_43 sn53_43 202000.000000
Rwneg53_44 in53_44 sn53_44 78000.000000
Rwneg53_45 in53_45 sn53_45 202000.000000
Rwneg53_46 in53_46 sn53_46 78000.000000
Rwneg53_47 in53_47 sn53_47 78000.000000
Rwneg53_48 in53_48 sn53_48 78000.000000
Rwneg53_49 in53_49 sn53_49 78000.000000
Rwneg53_50 in53_50 sn53_50 202000.000000
Rwneg53_51 in53_51 sn53_51 78000.000000
Rwneg53_52 in53_52 sn53_52 78000.000000
Rwneg53_53 in53_53 sn53_53 78000.000000
Rwneg53_54 in53_54 sn53_54 202000.000000
Rwneg53_55 in53_55 sn53_55 78000.000000
Rwneg53_56 in53_56 sn53_56 202000.000000
Rwneg53_57 in53_57 sn53_57 78000.000000
Rwneg53_58 in53_58 sn53_58 202000.000000
Rwneg53_59 in53_59 sn53_59 202000.000000
Rwneg53_60 in53_60 sn53_60 78000.000000
Rwneg53_61 in53_61 sn53_61 78000.000000
Rwneg53_62 in53_62 sn53_62 202000.000000
Rwneg53_63 in53_63 sn53_63 78000.000000
Rwneg53_64 in53_64 sn53_64 78000.000000
Rwneg53_65 in53_65 sn53_65 202000.000000
Rwneg53_66 in53_66 sn53_66 202000.000000
Rwneg53_67 in53_67 sn53_67 78000.000000
Rwneg53_68 in53_68 sn53_68 202000.000000
Rwneg53_69 in53_69 sn53_69 78000.000000
Rwneg53_70 in53_70 sn53_70 78000.000000
Rwneg53_71 in53_71 sn53_71 202000.000000
Rwneg53_72 in53_72 sn53_72 78000.000000
Rwneg53_73 in53_73 sn53_73 78000.000000
Rwneg53_74 in53_74 sn53_74 78000.000000
Rwneg53_75 in53_75 sn53_75 78000.000000
Rwneg53_76 in53_76 sn53_76 78000.000000
Rwneg53_77 in53_77 sn53_77 202000.000000
Rwneg53_78 in53_78 sn53_78 202000.000000
Rwneg53_79 in53_79 sn53_79 202000.000000
Rwneg53_80 in53_80 sn53_80 202000.000000
Rwneg53_81 in53_81 sn53_81 202000.000000
Rwneg53_82 in53_82 sn53_82 78000.000000
Rwneg53_83 in53_83 sn53_83 202000.000000
Rwneg53_84 in53_84 sn53_84 202000.000000
Rwneg54_1 in54_1 sn54_1 78000.000000
Rwneg54_2 in54_2 sn54_2 202000.000000
Rwneg54_3 in54_3 sn54_3 202000.000000
Rwneg54_4 in54_4 sn54_4 78000.000000
Rwneg54_5 in54_5 sn54_5 78000.000000
Rwneg54_6 in54_6 sn54_6 202000.000000
Rwneg54_7 in54_7 sn54_7 202000.000000
Rwneg54_8 in54_8 sn54_8 202000.000000
Rwneg54_9 in54_9 sn54_9 202000.000000
Rwneg54_10 in54_10 sn54_10 202000.000000
Rwneg54_11 in54_11 sn54_11 202000.000000
Rwneg54_12 in54_12 sn54_12 78000.000000
Rwneg54_13 in54_13 sn54_13 78000.000000
Rwneg54_14 in54_14 sn54_14 202000.000000
Rwneg54_15 in54_15 sn54_15 78000.000000
Rwneg54_16 in54_16 sn54_16 78000.000000
Rwneg54_17 in54_17 sn54_17 202000.000000
Rwneg54_18 in54_18 sn54_18 78000.000000
Rwneg54_19 in54_19 sn54_19 78000.000000
Rwneg54_20 in54_20 sn54_20 78000.000000
Rwneg54_21 in54_21 sn54_21 202000.000000
Rwneg54_22 in54_22 sn54_22 78000.000000
Rwneg54_23 in54_23 sn54_23 202000.000000
Rwneg54_24 in54_24 sn54_24 78000.000000
Rwneg54_25 in54_25 sn54_25 202000.000000
Rwneg54_26 in54_26 sn54_26 78000.000000
Rwneg54_27 in54_27 sn54_27 78000.000000
Rwneg54_28 in54_28 sn54_28 78000.000000
Rwneg54_29 in54_29 sn54_29 202000.000000
Rwneg54_30 in54_30 sn54_30 202000.000000
Rwneg54_31 in54_31 sn54_31 78000.000000
Rwneg54_32 in54_32 sn54_32 78000.000000
Rwneg54_33 in54_33 sn54_33 202000.000000
Rwneg54_34 in54_34 sn54_34 202000.000000
Rwneg54_35 in54_35 sn54_35 202000.000000
Rwneg54_36 in54_36 sn54_36 202000.000000
Rwneg54_37 in54_37 sn54_37 202000.000000
Rwneg54_38 in54_38 sn54_38 78000.000000
Rwneg54_39 in54_39 sn54_39 78000.000000
Rwneg54_40 in54_40 sn54_40 78000.000000
Rwneg54_41 in54_41 sn54_41 78000.000000
Rwneg54_42 in54_42 sn54_42 202000.000000
Rwneg54_43 in54_43 sn54_43 202000.000000
Rwneg54_44 in54_44 sn54_44 202000.000000
Rwneg54_45 in54_45 sn54_45 78000.000000
Rwneg54_46 in54_46 sn54_46 78000.000000
Rwneg54_47 in54_47 sn54_47 202000.000000
Rwneg54_48 in54_48 sn54_48 78000.000000
Rwneg54_49 in54_49 sn54_49 202000.000000
Rwneg54_50 in54_50 sn54_50 202000.000000
Rwneg54_51 in54_51 sn54_51 78000.000000
Rwneg54_52 in54_52 sn54_52 202000.000000
Rwneg54_53 in54_53 sn54_53 78000.000000
Rwneg54_54 in54_54 sn54_54 78000.000000
Rwneg54_55 in54_55 sn54_55 78000.000000
Rwneg54_56 in54_56 sn54_56 78000.000000
Rwneg54_57 in54_57 sn54_57 202000.000000
Rwneg54_58 in54_58 sn54_58 202000.000000
Rwneg54_59 in54_59 sn54_59 202000.000000
Rwneg54_60 in54_60 sn54_60 202000.000000
Rwneg54_61 in54_61 sn54_61 202000.000000
Rwneg54_62 in54_62 sn54_62 78000.000000
Rwneg54_63 in54_63 sn54_63 202000.000000
Rwneg54_64 in54_64 sn54_64 78000.000000
Rwneg54_65 in54_65 sn54_65 202000.000000
Rwneg54_66 in54_66 sn54_66 78000.000000
Rwneg54_67 in54_67 sn54_67 78000.000000
Rwneg54_68 in54_68 sn54_68 202000.000000
Rwneg54_69 in54_69 sn54_69 78000.000000
Rwneg54_70 in54_70 sn54_70 78000.000000
Rwneg54_71 in54_71 sn54_71 202000.000000
Rwneg54_72 in54_72 sn54_72 202000.000000
Rwneg54_73 in54_73 sn54_73 202000.000000
Rwneg54_74 in54_74 sn54_74 202000.000000
Rwneg54_75 in54_75 sn54_75 78000.000000
Rwneg54_76 in54_76 sn54_76 202000.000000
Rwneg54_77 in54_77 sn54_77 202000.000000
Rwneg54_78 in54_78 sn54_78 78000.000000
Rwneg54_79 in54_79 sn54_79 78000.000000
Rwneg54_80 in54_80 sn54_80 78000.000000
Rwneg54_81 in54_81 sn54_81 202000.000000
Rwneg54_82 in54_82 sn54_82 202000.000000
Rwneg54_83 in54_83 sn54_83 202000.000000
Rwneg54_84 in54_84 sn54_84 202000.000000
Rwneg55_1 in55_1 sn55_1 78000.000000
Rwneg55_2 in55_2 sn55_2 78000.000000
Rwneg55_3 in55_3 sn55_3 78000.000000
Rwneg55_4 in55_4 sn55_4 78000.000000
Rwneg55_5 in55_5 sn55_5 78000.000000
Rwneg55_6 in55_6 sn55_6 202000.000000
Rwneg55_7 in55_7 sn55_7 202000.000000
Rwneg55_8 in55_8 sn55_8 78000.000000
Rwneg55_9 in55_9 sn55_9 78000.000000
Rwneg55_10 in55_10 sn55_10 78000.000000
Rwneg55_11 in55_11 sn55_11 202000.000000
Rwneg55_12 in55_12 sn55_12 78000.000000
Rwneg55_13 in55_13 sn55_13 202000.000000
Rwneg55_14 in55_14 sn55_14 202000.000000
Rwneg55_15 in55_15 sn55_15 202000.000000
Rwneg55_16 in55_16 sn55_16 78000.000000
Rwneg55_17 in55_17 sn55_17 202000.000000
Rwneg55_18 in55_18 sn55_18 78000.000000
Rwneg55_19 in55_19 sn55_19 202000.000000
Rwneg55_20 in55_20 sn55_20 78000.000000
Rwneg55_21 in55_21 sn55_21 202000.000000
Rwneg55_22 in55_22 sn55_22 78000.000000
Rwneg55_23 in55_23 sn55_23 202000.000000
Rwneg55_24 in55_24 sn55_24 202000.000000
Rwneg55_25 in55_25 sn55_25 78000.000000
Rwneg55_26 in55_26 sn55_26 78000.000000
Rwneg55_27 in55_27 sn55_27 78000.000000
Rwneg55_28 in55_28 sn55_28 78000.000000
Rwneg55_29 in55_29 sn55_29 202000.000000
Rwneg55_30 in55_30 sn55_30 202000.000000
Rwneg55_31 in55_31 sn55_31 202000.000000
Rwneg55_32 in55_32 sn55_32 202000.000000
Rwneg55_33 in55_33 sn55_33 78000.000000
Rwneg55_34 in55_34 sn55_34 78000.000000
Rwneg55_35 in55_35 sn55_35 202000.000000
Rwneg55_36 in55_36 sn55_36 202000.000000
Rwneg55_37 in55_37 sn55_37 78000.000000
Rwneg55_38 in55_38 sn55_38 202000.000000
Rwneg55_39 in55_39 sn55_39 202000.000000
Rwneg55_40 in55_40 sn55_40 202000.000000
Rwneg55_41 in55_41 sn55_41 202000.000000
Rwneg55_42 in55_42 sn55_42 78000.000000
Rwneg55_43 in55_43 sn55_43 78000.000000
Rwneg55_44 in55_44 sn55_44 202000.000000
Rwneg55_45 in55_45 sn55_45 78000.000000
Rwneg55_46 in55_46 sn55_46 202000.000000
Rwneg55_47 in55_47 sn55_47 202000.000000
Rwneg55_48 in55_48 sn55_48 202000.000000
Rwneg55_49 in55_49 sn55_49 78000.000000
Rwneg55_50 in55_50 sn55_50 78000.000000
Rwneg55_51 in55_51 sn55_51 202000.000000
Rwneg55_52 in55_52 sn55_52 78000.000000
Rwneg55_53 in55_53 sn55_53 202000.000000
Rwneg55_54 in55_54 sn55_54 78000.000000
Rwneg55_55 in55_55 sn55_55 78000.000000
Rwneg55_56 in55_56 sn55_56 202000.000000
Rwneg55_57 in55_57 sn55_57 202000.000000
Rwneg55_58 in55_58 sn55_58 202000.000000
Rwneg55_59 in55_59 sn55_59 202000.000000
Rwneg55_60 in55_60 sn55_60 202000.000000
Rwneg55_61 in55_61 sn55_61 78000.000000
Rwneg55_62 in55_62 sn55_62 202000.000000
Rwneg55_63 in55_63 sn55_63 202000.000000
Rwneg55_64 in55_64 sn55_64 78000.000000
Rwneg55_65 in55_65 sn55_65 202000.000000
Rwneg55_66 in55_66 sn55_66 202000.000000
Rwneg55_67 in55_67 sn55_67 202000.000000
Rwneg55_68 in55_68 sn55_68 202000.000000
Rwneg55_69 in55_69 sn55_69 78000.000000
Rwneg55_70 in55_70 sn55_70 202000.000000
Rwneg55_71 in55_71 sn55_71 78000.000000
Rwneg55_72 in55_72 sn55_72 202000.000000
Rwneg55_73 in55_73 sn55_73 202000.000000
Rwneg55_74 in55_74 sn55_74 202000.000000
Rwneg55_75 in55_75 sn55_75 202000.000000
Rwneg55_76 in55_76 sn55_76 202000.000000
Rwneg55_77 in55_77 sn55_77 202000.000000
Rwneg55_78 in55_78 sn55_78 78000.000000
Rwneg55_79 in55_79 sn55_79 202000.000000
Rwneg55_80 in55_80 sn55_80 78000.000000
Rwneg55_81 in55_81 sn55_81 202000.000000
Rwneg55_82 in55_82 sn55_82 78000.000000
Rwneg55_83 in55_83 sn55_83 78000.000000
Rwneg55_84 in55_84 sn55_84 78000.000000
Rwneg56_1 in56_1 sn56_1 78000.000000
Rwneg56_2 in56_2 sn56_2 202000.000000
Rwneg56_3 in56_3 sn56_3 78000.000000
Rwneg56_4 in56_4 sn56_4 78000.000000
Rwneg56_5 in56_5 sn56_5 202000.000000
Rwneg56_6 in56_6 sn56_6 202000.000000
Rwneg56_7 in56_7 sn56_7 202000.000000
Rwneg56_8 in56_8 sn56_8 202000.000000
Rwneg56_9 in56_9 sn56_9 202000.000000
Rwneg56_10 in56_10 sn56_10 78000.000000
Rwneg56_11 in56_11 sn56_11 78000.000000
Rwneg56_12 in56_12 sn56_12 78000.000000
Rwneg56_13 in56_13 sn56_13 78000.000000
Rwneg56_14 in56_14 sn56_14 78000.000000
Rwneg56_15 in56_15 sn56_15 78000.000000
Rwneg56_16 in56_16 sn56_16 78000.000000
Rwneg56_17 in56_17 sn56_17 202000.000000
Rwneg56_18 in56_18 sn56_18 202000.000000
Rwneg56_19 in56_19 sn56_19 202000.000000
Rwneg56_20 in56_20 sn56_20 78000.000000
Rwneg56_21 in56_21 sn56_21 202000.000000
Rwneg56_22 in56_22 sn56_22 78000.000000
Rwneg56_23 in56_23 sn56_23 202000.000000
Rwneg56_24 in56_24 sn56_24 78000.000000
Rwneg56_25 in56_25 sn56_25 202000.000000
Rwneg56_26 in56_26 sn56_26 202000.000000
Rwneg56_27 in56_27 sn56_27 78000.000000
Rwneg56_28 in56_28 sn56_28 78000.000000
Rwneg56_29 in56_29 sn56_29 78000.000000
Rwneg56_30 in56_30 sn56_30 202000.000000
Rwneg56_31 in56_31 sn56_31 78000.000000
Rwneg56_32 in56_32 sn56_32 202000.000000
Rwneg56_33 in56_33 sn56_33 78000.000000
Rwneg56_34 in56_34 sn56_34 202000.000000
Rwneg56_35 in56_35 sn56_35 78000.000000
Rwneg56_36 in56_36 sn56_36 202000.000000
Rwneg56_37 in56_37 sn56_37 202000.000000
Rwneg56_38 in56_38 sn56_38 78000.000000
Rwneg56_39 in56_39 sn56_39 78000.000000
Rwneg56_40 in56_40 sn56_40 202000.000000
Rwneg56_41 in56_41 sn56_41 78000.000000
Rwneg56_42 in56_42 sn56_42 202000.000000
Rwneg56_43 in56_43 sn56_43 78000.000000
Rwneg56_44 in56_44 sn56_44 202000.000000
Rwneg56_45 in56_45 sn56_45 78000.000000
Rwneg56_46 in56_46 sn56_46 78000.000000
Rwneg56_47 in56_47 sn56_47 78000.000000
Rwneg56_48 in56_48 sn56_48 202000.000000
Rwneg56_49 in56_49 sn56_49 202000.000000
Rwneg56_50 in56_50 sn56_50 78000.000000
Rwneg56_51 in56_51 sn56_51 202000.000000
Rwneg56_52 in56_52 sn56_52 78000.000000
Rwneg56_53 in56_53 sn56_53 202000.000000
Rwneg56_54 in56_54 sn56_54 202000.000000
Rwneg56_55 in56_55 sn56_55 78000.000000
Rwneg56_56 in56_56 sn56_56 202000.000000
Rwneg56_57 in56_57 sn56_57 78000.000000
Rwneg56_58 in56_58 sn56_58 202000.000000
Rwneg56_59 in56_59 sn56_59 202000.000000
Rwneg56_60 in56_60 sn56_60 202000.000000
Rwneg56_61 in56_61 sn56_61 202000.000000
Rwneg56_62 in56_62 sn56_62 202000.000000
Rwneg56_63 in56_63 sn56_63 202000.000000
Rwneg56_64 in56_64 sn56_64 78000.000000
Rwneg56_65 in56_65 sn56_65 202000.000000
Rwneg56_66 in56_66 sn56_66 202000.000000
Rwneg56_67 in56_67 sn56_67 78000.000000
Rwneg56_68 in56_68 sn56_68 202000.000000
Rwneg56_69 in56_69 sn56_69 202000.000000
Rwneg56_70 in56_70 sn56_70 78000.000000
Rwneg56_71 in56_71 sn56_71 202000.000000
Rwneg56_72 in56_72 sn56_72 78000.000000
Rwneg56_73 in56_73 sn56_73 202000.000000
Rwneg56_74 in56_74 sn56_74 78000.000000
Rwneg56_75 in56_75 sn56_75 78000.000000
Rwneg56_76 in56_76 sn56_76 202000.000000
Rwneg56_77 in56_77 sn56_77 202000.000000
Rwneg56_78 in56_78 sn56_78 78000.000000
Rwneg56_79 in56_79 sn56_79 202000.000000
Rwneg56_80 in56_80 sn56_80 202000.000000
Rwneg56_81 in56_81 sn56_81 202000.000000
Rwneg56_82 in56_82 sn56_82 202000.000000
Rwneg56_83 in56_83 sn56_83 202000.000000
Rwneg56_84 in56_84 sn56_84 78000.000000
Rwneg57_1 in57_1 sn57_1 202000.000000
Rwneg57_2 in57_2 sn57_2 78000.000000
Rwneg57_3 in57_3 sn57_3 202000.000000
Rwneg57_4 in57_4 sn57_4 202000.000000
Rwneg57_5 in57_5 sn57_5 202000.000000
Rwneg57_6 in57_6 sn57_6 78000.000000
Rwneg57_7 in57_7 sn57_7 78000.000000
Rwneg57_8 in57_8 sn57_8 78000.000000
Rwneg57_9 in57_9 sn57_9 202000.000000
Rwneg57_10 in57_10 sn57_10 78000.000000
Rwneg57_11 in57_11 sn57_11 202000.000000
Rwneg57_12 in57_12 sn57_12 202000.000000
Rwneg57_13 in57_13 sn57_13 78000.000000
Rwneg57_14 in57_14 sn57_14 78000.000000
Rwneg57_15 in57_15 sn57_15 202000.000000
Rwneg57_16 in57_16 sn57_16 78000.000000
Rwneg57_17 in57_17 sn57_17 202000.000000
Rwneg57_18 in57_18 sn57_18 78000.000000
Rwneg57_19 in57_19 sn57_19 78000.000000
Rwneg57_20 in57_20 sn57_20 78000.000000
Rwneg57_21 in57_21 sn57_21 202000.000000
Rwneg57_22 in57_22 sn57_22 202000.000000
Rwneg57_23 in57_23 sn57_23 202000.000000
Rwneg57_24 in57_24 sn57_24 202000.000000
Rwneg57_25 in57_25 sn57_25 202000.000000
Rwneg57_26 in57_26 sn57_26 78000.000000
Rwneg57_27 in57_27 sn57_27 202000.000000
Rwneg57_28 in57_28 sn57_28 78000.000000
Rwneg57_29 in57_29 sn57_29 78000.000000
Rwneg57_30 in57_30 sn57_30 78000.000000
Rwneg57_31 in57_31 sn57_31 202000.000000
Rwneg57_32 in57_32 sn57_32 202000.000000
Rwneg57_33 in57_33 sn57_33 78000.000000
Rwneg57_34 in57_34 sn57_34 78000.000000
Rwneg57_35 in57_35 sn57_35 78000.000000
Rwneg57_36 in57_36 sn57_36 78000.000000
Rwneg57_37 in57_37 sn57_37 202000.000000
Rwneg57_38 in57_38 sn57_38 78000.000000
Rwneg57_39 in57_39 sn57_39 78000.000000
Rwneg57_40 in57_40 sn57_40 78000.000000
Rwneg57_41 in57_41 sn57_41 78000.000000
Rwneg57_42 in57_42 sn57_42 78000.000000
Rwneg57_43 in57_43 sn57_43 202000.000000
Rwneg57_44 in57_44 sn57_44 202000.000000
Rwneg57_45 in57_45 sn57_45 78000.000000
Rwneg57_46 in57_46 sn57_46 78000.000000
Rwneg57_47 in57_47 sn57_47 78000.000000
Rwneg57_48 in57_48 sn57_48 78000.000000
Rwneg57_49 in57_49 sn57_49 78000.000000
Rwneg57_50 in57_50 sn57_50 78000.000000
Rwneg57_51 in57_51 sn57_51 202000.000000
Rwneg57_52 in57_52 sn57_52 78000.000000
Rwneg57_53 in57_53 sn57_53 202000.000000
Rwneg57_54 in57_54 sn57_54 202000.000000
Rwneg57_55 in57_55 sn57_55 78000.000000
Rwneg57_56 in57_56 sn57_56 202000.000000
Rwneg57_57 in57_57 sn57_57 202000.000000
Rwneg57_58 in57_58 sn57_58 202000.000000
Rwneg57_59 in57_59 sn57_59 78000.000000
Rwneg57_60 in57_60 sn57_60 78000.000000
Rwneg57_61 in57_61 sn57_61 202000.000000
Rwneg57_62 in57_62 sn57_62 202000.000000
Rwneg57_63 in57_63 sn57_63 202000.000000
Rwneg57_64 in57_64 sn57_64 202000.000000
Rwneg57_65 in57_65 sn57_65 202000.000000
Rwneg57_66 in57_66 sn57_66 202000.000000
Rwneg57_67 in57_67 sn57_67 78000.000000
Rwneg57_68 in57_68 sn57_68 202000.000000
Rwneg57_69 in57_69 sn57_69 202000.000000
Rwneg57_70 in57_70 sn57_70 202000.000000
Rwneg57_71 in57_71 sn57_71 78000.000000
Rwneg57_72 in57_72 sn57_72 202000.000000
Rwneg57_73 in57_73 sn57_73 202000.000000
Rwneg57_74 in57_74 sn57_74 202000.000000
Rwneg57_75 in57_75 sn57_75 78000.000000
Rwneg57_76 in57_76 sn57_76 78000.000000
Rwneg57_77 in57_77 sn57_77 78000.000000
Rwneg57_78 in57_78 sn57_78 202000.000000
Rwneg57_79 in57_79 sn57_79 202000.000000
Rwneg57_80 in57_80 sn57_80 202000.000000
Rwneg57_81 in57_81 sn57_81 202000.000000
Rwneg57_82 in57_82 sn57_82 202000.000000
Rwneg57_83 in57_83 sn57_83 78000.000000
Rwneg57_84 in57_84 sn57_84 202000.000000
Rwneg58_1 in58_1 sn58_1 202000.000000
Rwneg58_2 in58_2 sn58_2 202000.000000
Rwneg58_3 in58_3 sn58_3 202000.000000
Rwneg58_4 in58_4 sn58_4 202000.000000
Rwneg58_5 in58_5 sn58_5 78000.000000
Rwneg58_6 in58_6 sn58_6 78000.000000
Rwneg58_7 in58_7 sn58_7 78000.000000
Rwneg58_8 in58_8 sn58_8 78000.000000
Rwneg58_9 in58_9 sn58_9 78000.000000
Rwneg58_10 in58_10 sn58_10 202000.000000
Rwneg58_11 in58_11 sn58_11 78000.000000
Rwneg58_12 in58_12 sn58_12 78000.000000
Rwneg58_13 in58_13 sn58_13 202000.000000
Rwneg58_14 in58_14 sn58_14 202000.000000
Rwneg58_15 in58_15 sn58_15 202000.000000
Rwneg58_16 in58_16 sn58_16 78000.000000
Rwneg58_17 in58_17 sn58_17 202000.000000
Rwneg58_18 in58_18 sn58_18 202000.000000
Rwneg58_19 in58_19 sn58_19 78000.000000
Rwneg58_20 in58_20 sn58_20 202000.000000
Rwneg58_21 in58_21 sn58_21 78000.000000
Rwneg58_22 in58_22 sn58_22 202000.000000
Rwneg58_23 in58_23 sn58_23 202000.000000
Rwneg58_24 in58_24 sn58_24 202000.000000
Rwneg58_25 in58_25 sn58_25 78000.000000
Rwneg58_26 in58_26 sn58_26 78000.000000
Rwneg58_27 in58_27 sn58_27 78000.000000
Rwneg58_28 in58_28 sn58_28 78000.000000
Rwneg58_29 in58_29 sn58_29 202000.000000
Rwneg58_30 in58_30 sn58_30 78000.000000
Rwneg58_31 in58_31 sn58_31 78000.000000
Rwneg58_32 in58_32 sn58_32 202000.000000
Rwneg58_33 in58_33 sn58_33 202000.000000
Rwneg58_34 in58_34 sn58_34 78000.000000
Rwneg58_35 in58_35 sn58_35 202000.000000
Rwneg58_36 in58_36 sn58_36 202000.000000
Rwneg58_37 in58_37 sn58_37 78000.000000
Rwneg58_38 in58_38 sn58_38 78000.000000
Rwneg58_39 in58_39 sn58_39 202000.000000
Rwneg58_40 in58_40 sn58_40 78000.000000
Rwneg58_41 in58_41 sn58_41 78000.000000
Rwneg58_42 in58_42 sn58_42 78000.000000
Rwneg58_43 in58_43 sn58_43 78000.000000
Rwneg58_44 in58_44 sn58_44 78000.000000
Rwneg58_45 in58_45 sn58_45 78000.000000
Rwneg58_46 in58_46 sn58_46 202000.000000
Rwneg58_47 in58_47 sn58_47 202000.000000
Rwneg58_48 in58_48 sn58_48 78000.000000
Rwneg58_49 in58_49 sn58_49 202000.000000
Rwneg58_50 in58_50 sn58_50 202000.000000
Rwneg58_51 in58_51 sn58_51 78000.000000
Rwneg58_52 in58_52 sn58_52 202000.000000
Rwneg58_53 in58_53 sn58_53 202000.000000
Rwneg58_54 in58_54 sn58_54 202000.000000
Rwneg58_55 in58_55 sn58_55 202000.000000
Rwneg58_56 in58_56 sn58_56 78000.000000
Rwneg58_57 in58_57 sn58_57 202000.000000
Rwneg58_58 in58_58 sn58_58 78000.000000
Rwneg58_59 in58_59 sn58_59 78000.000000
Rwneg58_60 in58_60 sn58_60 202000.000000
Rwneg58_61 in58_61 sn58_61 78000.000000
Rwneg58_62 in58_62 sn58_62 202000.000000
Rwneg58_63 in58_63 sn58_63 78000.000000
Rwneg58_64 in58_64 sn58_64 202000.000000
Rwneg58_65 in58_65 sn58_65 78000.000000
Rwneg58_66 in58_66 sn58_66 78000.000000
Rwneg58_67 in58_67 sn58_67 202000.000000
Rwneg58_68 in58_68 sn58_68 78000.000000
Rwneg58_69 in58_69 sn58_69 78000.000000
Rwneg58_70 in58_70 sn58_70 78000.000000
Rwneg58_71 in58_71 sn58_71 78000.000000
Rwneg58_72 in58_72 sn58_72 78000.000000
Rwneg58_73 in58_73 sn58_73 78000.000000
Rwneg58_74 in58_74 sn58_74 202000.000000
Rwneg58_75 in58_75 sn58_75 202000.000000
Rwneg58_76 in58_76 sn58_76 78000.000000
Rwneg58_77 in58_77 sn58_77 78000.000000
Rwneg58_78 in58_78 sn58_78 202000.000000
Rwneg58_79 in58_79 sn58_79 202000.000000
Rwneg58_80 in58_80 sn58_80 78000.000000
Rwneg58_81 in58_81 sn58_81 202000.000000
Rwneg58_82 in58_82 sn58_82 78000.000000
Rwneg58_83 in58_83 sn58_83 202000.000000
Rwneg58_84 in58_84 sn58_84 202000.000000
Rwneg59_1 in59_1 sn59_1 202000.000000
Rwneg59_2 in59_2 sn59_2 78000.000000
Rwneg59_3 in59_3 sn59_3 78000.000000
Rwneg59_4 in59_4 sn59_4 78000.000000
Rwneg59_5 in59_5 sn59_5 78000.000000
Rwneg59_6 in59_6 sn59_6 202000.000000
Rwneg59_7 in59_7 sn59_7 202000.000000
Rwneg59_8 in59_8 sn59_8 78000.000000
Rwneg59_9 in59_9 sn59_9 78000.000000
Rwneg59_10 in59_10 sn59_10 202000.000000
Rwneg59_11 in59_11 sn59_11 202000.000000
Rwneg59_12 in59_12 sn59_12 202000.000000
Rwneg59_13 in59_13 sn59_13 78000.000000
Rwneg59_14 in59_14 sn59_14 78000.000000
Rwneg59_15 in59_15 sn59_15 78000.000000
Rwneg59_16 in59_16 sn59_16 202000.000000
Rwneg59_17 in59_17 sn59_17 202000.000000
Rwneg59_18 in59_18 sn59_18 202000.000000
Rwneg59_19 in59_19 sn59_19 78000.000000
Rwneg59_20 in59_20 sn59_20 78000.000000
Rwneg59_21 in59_21 sn59_21 202000.000000
Rwneg59_22 in59_22 sn59_22 202000.000000
Rwneg59_23 in59_23 sn59_23 202000.000000
Rwneg59_24 in59_24 sn59_24 202000.000000
Rwneg59_25 in59_25 sn59_25 202000.000000
Rwneg59_26 in59_26 sn59_26 78000.000000
Rwneg59_27 in59_27 sn59_27 78000.000000
Rwneg59_28 in59_28 sn59_28 202000.000000
Rwneg59_29 in59_29 sn59_29 202000.000000
Rwneg59_30 in59_30 sn59_30 202000.000000
Rwneg59_31 in59_31 sn59_31 78000.000000
Rwneg59_32 in59_32 sn59_32 202000.000000
Rwneg59_33 in59_33 sn59_33 78000.000000
Rwneg59_34 in59_34 sn59_34 202000.000000
Rwneg59_35 in59_35 sn59_35 202000.000000
Rwneg59_36 in59_36 sn59_36 202000.000000
Rwneg59_37 in59_37 sn59_37 202000.000000
Rwneg59_38 in59_38 sn59_38 78000.000000
Rwneg59_39 in59_39 sn59_39 202000.000000
Rwneg59_40 in59_40 sn59_40 202000.000000
Rwneg59_41 in59_41 sn59_41 202000.000000
Rwneg59_42 in59_42 sn59_42 78000.000000
Rwneg59_43 in59_43 sn59_43 78000.000000
Rwneg59_44 in59_44 sn59_44 78000.000000
Rwneg59_45 in59_45 sn59_45 78000.000000
Rwneg59_46 in59_46 sn59_46 202000.000000
Rwneg59_47 in59_47 sn59_47 202000.000000
Rwneg59_48 in59_48 sn59_48 202000.000000
Rwneg59_49 in59_49 sn59_49 78000.000000
Rwneg59_50 in59_50 sn59_50 78000.000000
Rwneg59_51 in59_51 sn59_51 202000.000000
Rwneg59_52 in59_52 sn59_52 78000.000000
Rwneg59_53 in59_53 sn59_53 202000.000000
Rwneg59_54 in59_54 sn59_54 78000.000000
Rwneg59_55 in59_55 sn59_55 78000.000000
Rwneg59_56 in59_56 sn59_56 78000.000000
Rwneg59_57 in59_57 sn59_57 78000.000000
Rwneg59_58 in59_58 sn59_58 202000.000000
Rwneg59_59 in59_59 sn59_59 202000.000000
Rwneg59_60 in59_60 sn59_60 78000.000000
Rwneg59_61 in59_61 sn59_61 78000.000000
Rwneg59_62 in59_62 sn59_62 202000.000000
Rwneg59_63 in59_63 sn59_63 78000.000000
Rwneg59_64 in59_64 sn59_64 202000.000000
Rwneg59_65 in59_65 sn59_65 202000.000000
Rwneg59_66 in59_66 sn59_66 78000.000000
Rwneg59_67 in59_67 sn59_67 202000.000000
Rwneg59_68 in59_68 sn59_68 202000.000000
Rwneg59_69 in59_69 sn59_69 78000.000000
Rwneg59_70 in59_70 sn59_70 202000.000000
Rwneg59_71 in59_71 sn59_71 78000.000000
Rwneg59_72 in59_72 sn59_72 202000.000000
Rwneg59_73 in59_73 sn59_73 202000.000000
Rwneg59_74 in59_74 sn59_74 202000.000000
Rwneg59_75 in59_75 sn59_75 202000.000000
Rwneg59_76 in59_76 sn59_76 78000.000000
Rwneg59_77 in59_77 sn59_77 202000.000000
Rwneg59_78 in59_78 sn59_78 78000.000000
Rwneg59_79 in59_79 sn59_79 202000.000000
Rwneg59_80 in59_80 sn59_80 202000.000000
Rwneg59_81 in59_81 sn59_81 202000.000000
Rwneg59_82 in59_82 sn59_82 202000.000000
Rwneg59_83 in59_83 sn59_83 78000.000000
Rwneg59_84 in59_84 sn59_84 202000.000000
Rwneg60_1 in60_1 sn60_1 202000.000000
Rwneg60_2 in60_2 sn60_2 202000.000000
Rwneg60_3 in60_3 sn60_3 202000.000000
Rwneg60_4 in60_4 sn60_4 202000.000000
Rwneg60_5 in60_5 sn60_5 78000.000000
Rwneg60_6 in60_6 sn60_6 78000.000000
Rwneg60_7 in60_7 sn60_7 202000.000000
Rwneg60_8 in60_8 sn60_8 202000.000000
Rwneg60_9 in60_9 sn60_9 78000.000000
Rwneg60_10 in60_10 sn60_10 202000.000000
Rwneg60_11 in60_11 sn60_11 202000.000000
Rwneg60_12 in60_12 sn60_12 78000.000000
Rwneg60_13 in60_13 sn60_13 78000.000000
Rwneg60_14 in60_14 sn60_14 78000.000000
Rwneg60_15 in60_15 sn60_15 78000.000000
Rwneg60_16 in60_16 sn60_16 202000.000000
Rwneg60_17 in60_17 sn60_17 78000.000000
Rwneg60_18 in60_18 sn60_18 78000.000000
Rwneg60_19 in60_19 sn60_19 78000.000000
Rwneg60_20 in60_20 sn60_20 202000.000000
Rwneg60_21 in60_21 sn60_21 202000.000000
Rwneg60_22 in60_22 sn60_22 78000.000000
Rwneg60_23 in60_23 sn60_23 202000.000000
Rwneg60_24 in60_24 sn60_24 202000.000000
Rwneg60_25 in60_25 sn60_25 78000.000000
Rwneg60_26 in60_26 sn60_26 202000.000000
Rwneg60_27 in60_27 sn60_27 202000.000000
Rwneg60_28 in60_28 sn60_28 202000.000000
Rwneg60_29 in60_29 sn60_29 202000.000000
Rwneg60_30 in60_30 sn60_30 78000.000000
Rwneg60_31 in60_31 sn60_31 78000.000000
Rwneg60_32 in60_32 sn60_32 78000.000000
Rwneg60_33 in60_33 sn60_33 202000.000000
Rwneg60_34 in60_34 sn60_34 78000.000000
Rwneg60_35 in60_35 sn60_35 202000.000000
Rwneg60_36 in60_36 sn60_36 78000.000000
Rwneg60_37 in60_37 sn60_37 202000.000000
Rwneg60_38 in60_38 sn60_38 78000.000000
Rwneg60_39 in60_39 sn60_39 78000.000000
Rwneg60_40 in60_40 sn60_40 78000.000000
Rwneg60_41 in60_41 sn60_41 78000.000000
Rwneg60_42 in60_42 sn60_42 202000.000000
Rwneg60_43 in60_43 sn60_43 78000.000000
Rwneg60_44 in60_44 sn60_44 202000.000000
Rwneg60_45 in60_45 sn60_45 78000.000000
Rwneg60_46 in60_46 sn60_46 202000.000000
Rwneg60_47 in60_47 sn60_47 78000.000000
Rwneg60_48 in60_48 sn60_48 202000.000000
Rwneg60_49 in60_49 sn60_49 202000.000000
Rwneg60_50 in60_50 sn60_50 78000.000000
Rwneg60_51 in60_51 sn60_51 202000.000000
Rwneg60_52 in60_52 sn60_52 202000.000000
Rwneg60_53 in60_53 sn60_53 78000.000000
Rwneg60_54 in60_54 sn60_54 202000.000000
Rwneg60_55 in60_55 sn60_55 202000.000000
Rwneg60_56 in60_56 sn60_56 78000.000000
Rwneg60_57 in60_57 sn60_57 202000.000000
Rwneg60_58 in60_58 sn60_58 202000.000000
Rwneg60_59 in60_59 sn60_59 78000.000000
Rwneg60_60 in60_60 sn60_60 202000.000000
Rwneg60_61 in60_61 sn60_61 78000.000000
Rwneg60_62 in60_62 sn60_62 202000.000000
Rwneg60_63 in60_63 sn60_63 78000.000000
Rwneg60_64 in60_64 sn60_64 78000.000000
Rwneg60_65 in60_65 sn60_65 202000.000000
Rwneg60_66 in60_66 sn60_66 202000.000000
Rwneg60_67 in60_67 sn60_67 78000.000000
Rwneg60_68 in60_68 sn60_68 78000.000000
Rwneg60_69 in60_69 sn60_69 202000.000000
Rwneg60_70 in60_70 sn60_70 202000.000000
Rwneg60_71 in60_71 sn60_71 78000.000000
Rwneg60_72 in60_72 sn60_72 78000.000000
Rwneg60_73 in60_73 sn60_73 78000.000000
Rwneg60_74 in60_74 sn60_74 78000.000000
Rwneg60_75 in60_75 sn60_75 78000.000000
Rwneg60_76 in60_76 sn60_76 202000.000000
Rwneg60_77 in60_77 sn60_77 78000.000000
Rwneg60_78 in60_78 sn60_78 78000.000000
Rwneg60_79 in60_79 sn60_79 78000.000000
Rwneg60_80 in60_80 sn60_80 78000.000000
Rwneg60_81 in60_81 sn60_81 202000.000000
Rwneg60_82 in60_82 sn60_82 202000.000000
Rwneg60_83 in60_83 sn60_83 78000.000000
Rwneg60_84 in60_84 sn60_84 202000.000000
Rwneg61_1 in61_1 sn61_1 202000.000000
Rwneg61_2 in61_2 sn61_2 78000.000000
Rwneg61_3 in61_3 sn61_3 202000.000000
Rwneg61_4 in61_4 sn61_4 202000.000000
Rwneg61_5 in61_5 sn61_5 202000.000000
Rwneg61_6 in61_6 sn61_6 202000.000000
Rwneg61_7 in61_7 sn61_7 202000.000000
Rwneg61_8 in61_8 sn61_8 78000.000000
Rwneg61_9 in61_9 sn61_9 202000.000000
Rwneg61_10 in61_10 sn61_10 202000.000000
Rwneg61_11 in61_11 sn61_11 78000.000000
Rwneg61_12 in61_12 sn61_12 202000.000000
Rwneg61_13 in61_13 sn61_13 202000.000000
Rwneg61_14 in61_14 sn61_14 202000.000000
Rwneg61_15 in61_15 sn61_15 202000.000000
Rwneg61_16 in61_16 sn61_16 78000.000000
Rwneg61_17 in61_17 sn61_17 202000.000000
Rwneg61_18 in61_18 sn61_18 202000.000000
Rwneg61_19 in61_19 sn61_19 78000.000000
Rwneg61_20 in61_20 sn61_20 78000.000000
Rwneg61_21 in61_21 sn61_21 202000.000000
Rwneg61_22 in61_22 sn61_22 202000.000000
Rwneg61_23 in61_23 sn61_23 78000.000000
Rwneg61_24 in61_24 sn61_24 202000.000000
Rwneg61_25 in61_25 sn61_25 202000.000000
Rwneg61_26 in61_26 sn61_26 78000.000000
Rwneg61_27 in61_27 sn61_27 202000.000000
Rwneg61_28 in61_28 sn61_28 78000.000000
Rwneg61_29 in61_29 sn61_29 202000.000000
Rwneg61_30 in61_30 sn61_30 202000.000000
Rwneg61_31 in61_31 sn61_31 202000.000000
Rwneg61_32 in61_32 sn61_32 78000.000000
Rwneg61_33 in61_33 sn61_33 78000.000000
Rwneg61_34 in61_34 sn61_34 78000.000000
Rwneg61_35 in61_35 sn61_35 78000.000000
Rwneg61_36 in61_36 sn61_36 202000.000000
Rwneg61_37 in61_37 sn61_37 78000.000000
Rwneg61_38 in61_38 sn61_38 78000.000000
Rwneg61_39 in61_39 sn61_39 78000.000000
Rwneg61_40 in61_40 sn61_40 78000.000000
Rwneg61_41 in61_41 sn61_41 202000.000000
Rwneg61_42 in61_42 sn61_42 78000.000000
Rwneg61_43 in61_43 sn61_43 202000.000000
Rwneg61_44 in61_44 sn61_44 202000.000000
Rwneg61_45 in61_45 sn61_45 78000.000000
Rwneg61_46 in61_46 sn61_46 78000.000000
Rwneg61_47 in61_47 sn61_47 202000.000000
Rwneg61_48 in61_48 sn61_48 78000.000000
Rwneg61_49 in61_49 sn61_49 78000.000000
Rwneg61_50 in61_50 sn61_50 202000.000000
Rwneg61_51 in61_51 sn61_51 78000.000000
Rwneg61_52 in61_52 sn61_52 202000.000000
Rwneg61_53 in61_53 sn61_53 78000.000000
Rwneg61_54 in61_54 sn61_54 78000.000000
Rwneg61_55 in61_55 sn61_55 78000.000000
Rwneg61_56 in61_56 sn61_56 202000.000000
Rwneg61_57 in61_57 sn61_57 202000.000000
Rwneg61_58 in61_58 sn61_58 202000.000000
Rwneg61_59 in61_59 sn61_59 202000.000000
Rwneg61_60 in61_60 sn61_60 202000.000000
Rwneg61_61 in61_61 sn61_61 202000.000000
Rwneg61_62 in61_62 sn61_62 202000.000000
Rwneg61_63 in61_63 sn61_63 202000.000000
Rwneg61_64 in61_64 sn61_64 202000.000000
Rwneg61_65 in61_65 sn61_65 78000.000000
Rwneg61_66 in61_66 sn61_66 78000.000000
Rwneg61_67 in61_67 sn61_67 202000.000000
Rwneg61_68 in61_68 sn61_68 202000.000000
Rwneg61_69 in61_69 sn61_69 202000.000000
Rwneg61_70 in61_70 sn61_70 78000.000000
Rwneg61_71 in61_71 sn61_71 202000.000000
Rwneg61_72 in61_72 sn61_72 202000.000000
Rwneg61_73 in61_73 sn61_73 78000.000000
Rwneg61_74 in61_74 sn61_74 202000.000000
Rwneg61_75 in61_75 sn61_75 78000.000000
Rwneg61_76 in61_76 sn61_76 202000.000000
Rwneg61_77 in61_77 sn61_77 78000.000000
Rwneg61_78 in61_78 sn61_78 202000.000000
Rwneg61_79 in61_79 sn61_79 78000.000000
Rwneg61_80 in61_80 sn61_80 78000.000000
Rwneg61_81 in61_81 sn61_81 202000.000000
Rwneg61_82 in61_82 sn61_82 202000.000000
Rwneg61_83 in61_83 sn61_83 202000.000000
Rwneg61_84 in61_84 sn61_84 78000.000000
Rwneg62_1 in62_1 sn62_1 202000.000000
Rwneg62_2 in62_2 sn62_2 78000.000000
Rwneg62_3 in62_3 sn62_3 78000.000000
Rwneg62_4 in62_4 sn62_4 78000.000000
Rwneg62_5 in62_5 sn62_5 78000.000000
Rwneg62_6 in62_6 sn62_6 202000.000000
Rwneg62_7 in62_7 sn62_7 78000.000000
Rwneg62_8 in62_8 sn62_8 78000.000000
Rwneg62_9 in62_9 sn62_9 78000.000000
Rwneg62_10 in62_10 sn62_10 202000.000000
Rwneg62_11 in62_11 sn62_11 202000.000000
Rwneg62_12 in62_12 sn62_12 202000.000000
Rwneg62_13 in62_13 sn62_13 202000.000000
Rwneg62_14 in62_14 sn62_14 78000.000000
Rwneg62_15 in62_15 sn62_15 78000.000000
Rwneg62_16 in62_16 sn62_16 78000.000000
Rwneg62_17 in62_17 sn62_17 202000.000000
Rwneg62_18 in62_18 sn62_18 202000.000000
Rwneg62_19 in62_19 sn62_19 202000.000000
Rwneg62_20 in62_20 sn62_20 202000.000000
Rwneg62_21 in62_21 sn62_21 78000.000000
Rwneg62_22 in62_22 sn62_22 202000.000000
Rwneg62_23 in62_23 sn62_23 202000.000000
Rwneg62_24 in62_24 sn62_24 78000.000000
Rwneg62_25 in62_25 sn62_25 202000.000000
Rwneg62_26 in62_26 sn62_26 202000.000000
Rwneg62_27 in62_27 sn62_27 202000.000000
Rwneg62_28 in62_28 sn62_28 202000.000000
Rwneg62_29 in62_29 sn62_29 78000.000000
Rwneg62_30 in62_30 sn62_30 202000.000000
Rwneg62_31 in62_31 sn62_31 202000.000000
Rwneg62_32 in62_32 sn62_32 202000.000000
Rwneg62_33 in62_33 sn62_33 202000.000000
Rwneg62_34 in62_34 sn62_34 78000.000000
Rwneg62_35 in62_35 sn62_35 78000.000000
Rwneg62_36 in62_36 sn62_36 78000.000000
Rwneg62_37 in62_37 sn62_37 202000.000000
Rwneg62_38 in62_38 sn62_38 78000.000000
Rwneg62_39 in62_39 sn62_39 78000.000000
Rwneg62_40 in62_40 sn62_40 202000.000000
Rwneg62_41 in62_41 sn62_41 78000.000000
Rwneg62_42 in62_42 sn62_42 78000.000000
Rwneg62_43 in62_43 sn62_43 78000.000000
Rwneg62_44 in62_44 sn62_44 78000.000000
Rwneg62_45 in62_45 sn62_45 202000.000000
Rwneg62_46 in62_46 sn62_46 78000.000000
Rwneg62_47 in62_47 sn62_47 78000.000000
Rwneg62_48 in62_48 sn62_48 202000.000000
Rwneg62_49 in62_49 sn62_49 78000.000000
Rwneg62_50 in62_50 sn62_50 78000.000000
Rwneg62_51 in62_51 sn62_51 202000.000000
Rwneg62_52 in62_52 sn62_52 78000.000000
Rwneg62_53 in62_53 sn62_53 78000.000000
Rwneg62_54 in62_54 sn62_54 202000.000000
Rwneg62_55 in62_55 sn62_55 202000.000000
Rwneg62_56 in62_56 sn62_56 202000.000000
Rwneg62_57 in62_57 sn62_57 78000.000000
Rwneg62_58 in62_58 sn62_58 202000.000000
Rwneg62_59 in62_59 sn62_59 78000.000000
Rwneg62_60 in62_60 sn62_60 78000.000000
Rwneg62_61 in62_61 sn62_61 202000.000000
Rwneg62_62 in62_62 sn62_62 202000.000000
Rwneg62_63 in62_63 sn62_63 202000.000000
Rwneg62_64 in62_64 sn62_64 202000.000000
Rwneg62_65 in62_65 sn62_65 78000.000000
Rwneg62_66 in62_66 sn62_66 202000.000000
Rwneg62_67 in62_67 sn62_67 202000.000000
Rwneg62_68 in62_68 sn62_68 78000.000000
Rwneg62_69 in62_69 sn62_69 202000.000000
Rwneg62_70 in62_70 sn62_70 202000.000000
Rwneg62_71 in62_71 sn62_71 202000.000000
Rwneg62_72 in62_72 sn62_72 78000.000000
Rwneg62_73 in62_73 sn62_73 202000.000000
Rwneg62_74 in62_74 sn62_74 78000.000000
Rwneg62_75 in62_75 sn62_75 202000.000000
Rwneg62_76 in62_76 sn62_76 78000.000000
Rwneg62_77 in62_77 sn62_77 202000.000000
Rwneg62_78 in62_78 sn62_78 78000.000000
Rwneg62_79 in62_79 sn62_79 202000.000000
Rwneg62_80 in62_80 sn62_80 202000.000000
Rwneg62_81 in62_81 sn62_81 202000.000000
Rwneg62_82 in62_82 sn62_82 202000.000000
Rwneg62_83 in62_83 sn62_83 202000.000000
Rwneg62_84 in62_84 sn62_84 202000.000000
Rwneg63_1 in63_1 sn63_1 78000.000000
Rwneg63_2 in63_2 sn63_2 78000.000000
Rwneg63_3 in63_3 sn63_3 78000.000000
Rwneg63_4 in63_4 sn63_4 78000.000000
Rwneg63_5 in63_5 sn63_5 78000.000000
Rwneg63_6 in63_6 sn63_6 202000.000000
Rwneg63_7 in63_7 sn63_7 202000.000000
Rwneg63_8 in63_8 sn63_8 78000.000000
Rwneg63_9 in63_9 sn63_9 78000.000000
Rwneg63_10 in63_10 sn63_10 202000.000000
Rwneg63_11 in63_11 sn63_11 78000.000000
Rwneg63_12 in63_12 sn63_12 202000.000000
Rwneg63_13 in63_13 sn63_13 78000.000000
Rwneg63_14 in63_14 sn63_14 202000.000000
Rwneg63_15 in63_15 sn63_15 202000.000000
Rwneg63_16 in63_16 sn63_16 202000.000000
Rwneg63_17 in63_17 sn63_17 78000.000000
Rwneg63_18 in63_18 sn63_18 78000.000000
Rwneg63_19 in63_19 sn63_19 202000.000000
Rwneg63_20 in63_20 sn63_20 202000.000000
Rwneg63_21 in63_21 sn63_21 202000.000000
Rwneg63_22 in63_22 sn63_22 78000.000000
Rwneg63_23 in63_23 sn63_23 78000.000000
Rwneg63_24 in63_24 sn63_24 202000.000000
Rwneg63_25 in63_25 sn63_25 202000.000000
Rwneg63_26 in63_26 sn63_26 202000.000000
Rwneg63_27 in63_27 sn63_27 202000.000000
Rwneg63_28 in63_28 sn63_28 202000.000000
Rwneg63_29 in63_29 sn63_29 202000.000000
Rwneg63_30 in63_30 sn63_30 202000.000000
Rwneg63_31 in63_31 sn63_31 78000.000000
Rwneg63_32 in63_32 sn63_32 202000.000000
Rwneg63_33 in63_33 sn63_33 78000.000000
Rwneg63_34 in63_34 sn63_34 202000.000000
Rwneg63_35 in63_35 sn63_35 78000.000000
Rwneg63_36 in63_36 sn63_36 202000.000000
Rwneg63_37 in63_37 sn63_37 202000.000000
Rwneg63_38 in63_38 sn63_38 202000.000000
Rwneg63_39 in63_39 sn63_39 202000.000000
Rwneg63_40 in63_40 sn63_40 202000.000000
Rwneg63_41 in63_41 sn63_41 78000.000000
Rwneg63_42 in63_42 sn63_42 78000.000000
Rwneg63_43 in63_43 sn63_43 202000.000000
Rwneg63_44 in63_44 sn63_44 202000.000000
Rwneg63_45 in63_45 sn63_45 202000.000000
Rwneg63_46 in63_46 sn63_46 202000.000000
Rwneg63_47 in63_47 sn63_47 202000.000000
Rwneg63_48 in63_48 sn63_48 202000.000000
Rwneg63_49 in63_49 sn63_49 202000.000000
Rwneg63_50 in63_50 sn63_50 202000.000000
Rwneg63_51 in63_51 sn63_51 202000.000000
Rwneg63_52 in63_52 sn63_52 202000.000000
Rwneg63_53 in63_53 sn63_53 78000.000000
Rwneg63_54 in63_54 sn63_54 78000.000000
Rwneg63_55 in63_55 sn63_55 78000.000000
Rwneg63_56 in63_56 sn63_56 78000.000000
Rwneg63_57 in63_57 sn63_57 78000.000000
Rwneg63_58 in63_58 sn63_58 78000.000000
Rwneg63_59 in63_59 sn63_59 78000.000000
Rwneg63_60 in63_60 sn63_60 202000.000000
Rwneg63_61 in63_61 sn63_61 78000.000000
Rwneg63_62 in63_62 sn63_62 78000.000000
Rwneg63_63 in63_63 sn63_63 202000.000000
Rwneg63_64 in63_64 sn63_64 78000.000000
Rwneg63_65 in63_65 sn63_65 78000.000000
Rwneg63_66 in63_66 sn63_66 202000.000000
Rwneg63_67 in63_67 sn63_67 202000.000000
Rwneg63_68 in63_68 sn63_68 202000.000000
Rwneg63_69 in63_69 sn63_69 78000.000000
Rwneg63_70 in63_70 sn63_70 202000.000000
Rwneg63_71 in63_71 sn63_71 78000.000000
Rwneg63_72 in63_72 sn63_72 202000.000000
Rwneg63_73 in63_73 sn63_73 78000.000000
Rwneg63_74 in63_74 sn63_74 78000.000000
Rwneg63_75 in63_75 sn63_75 78000.000000
Rwneg63_76 in63_76 sn63_76 202000.000000
Rwneg63_77 in63_77 sn63_77 78000.000000
Rwneg63_78 in63_78 sn63_78 78000.000000
Rwneg63_79 in63_79 sn63_79 202000.000000
Rwneg63_80 in63_80 sn63_80 78000.000000
Rwneg63_81 in63_81 sn63_81 78000.000000
Rwneg63_82 in63_82 sn63_82 202000.000000
Rwneg63_83 in63_83 sn63_83 78000.000000
Rwneg63_84 in63_84 sn63_84 78000.000000
Rwneg64_1 in64_1 sn64_1 202000.000000
Rwneg64_2 in64_2 sn64_2 202000.000000
Rwneg64_3 in64_3 sn64_3 202000.000000
Rwneg64_4 in64_4 sn64_4 202000.000000
Rwneg64_5 in64_5 sn64_5 78000.000000
Rwneg64_6 in64_6 sn64_6 202000.000000
Rwneg64_7 in64_7 sn64_7 202000.000000
Rwneg64_8 in64_8 sn64_8 202000.000000
Rwneg64_9 in64_9 sn64_9 202000.000000
Rwneg64_10 in64_10 sn64_10 202000.000000
Rwneg64_11 in64_11 sn64_11 78000.000000
Rwneg64_12 in64_12 sn64_12 78000.000000
Rwneg64_13 in64_13 sn64_13 78000.000000
Rwneg64_14 in64_14 sn64_14 202000.000000
Rwneg64_15 in64_15 sn64_15 202000.000000
Rwneg64_16 in64_16 sn64_16 202000.000000
Rwneg64_17 in64_17 sn64_17 202000.000000
Rwneg64_18 in64_18 sn64_18 78000.000000
Rwneg64_19 in64_19 sn64_19 78000.000000
Rwneg64_20 in64_20 sn64_20 78000.000000
Rwneg64_21 in64_21 sn64_21 202000.000000
Rwneg64_22 in64_22 sn64_22 202000.000000
Rwneg64_23 in64_23 sn64_23 78000.000000
Rwneg64_24 in64_24 sn64_24 78000.000000
Rwneg64_25 in64_25 sn64_25 78000.000000
Rwneg64_26 in64_26 sn64_26 202000.000000
Rwneg64_27 in64_27 sn64_27 202000.000000
Rwneg64_28 in64_28 sn64_28 78000.000000
Rwneg64_29 in64_29 sn64_29 78000.000000
Rwneg64_30 in64_30 sn64_30 202000.000000
Rwneg64_31 in64_31 sn64_31 202000.000000
Rwneg64_32 in64_32 sn64_32 202000.000000
Rwneg64_33 in64_33 sn64_33 202000.000000
Rwneg64_34 in64_34 sn64_34 78000.000000
Rwneg64_35 in64_35 sn64_35 202000.000000
Rwneg64_36 in64_36 sn64_36 78000.000000
Rwneg64_37 in64_37 sn64_37 78000.000000
Rwneg64_38 in64_38 sn64_38 202000.000000
Rwneg64_39 in64_39 sn64_39 78000.000000
Rwneg64_40 in64_40 sn64_40 78000.000000
Rwneg64_41 in64_41 sn64_41 202000.000000
Rwneg64_42 in64_42 sn64_42 202000.000000
Rwneg64_43 in64_43 sn64_43 78000.000000
Rwneg64_44 in64_44 sn64_44 202000.000000
Rwneg64_45 in64_45 sn64_45 202000.000000
Rwneg64_46 in64_46 sn64_46 202000.000000
Rwneg64_47 in64_47 sn64_47 202000.000000
Rwneg64_48 in64_48 sn64_48 202000.000000
Rwneg64_49 in64_49 sn64_49 78000.000000
Rwneg64_50 in64_50 sn64_50 202000.000000
Rwneg64_51 in64_51 sn64_51 202000.000000
Rwneg64_52 in64_52 sn64_52 202000.000000
Rwneg64_53 in64_53 sn64_53 78000.000000
Rwneg64_54 in64_54 sn64_54 78000.000000
Rwneg64_55 in64_55 sn64_55 78000.000000
Rwneg64_56 in64_56 sn64_56 78000.000000
Rwneg64_57 in64_57 sn64_57 202000.000000
Rwneg64_58 in64_58 sn64_58 202000.000000
Rwneg64_59 in64_59 sn64_59 78000.000000
Rwneg64_60 in64_60 sn64_60 202000.000000
Rwneg64_61 in64_61 sn64_61 202000.000000
Rwneg64_62 in64_62 sn64_62 78000.000000
Rwneg64_63 in64_63 sn64_63 78000.000000
Rwneg64_64 in64_64 sn64_64 202000.000000
Rwneg64_65 in64_65 sn64_65 78000.000000
Rwneg64_66 in64_66 sn64_66 78000.000000
Rwneg64_67 in64_67 sn64_67 202000.000000
Rwneg64_68 in64_68 sn64_68 78000.000000
Rwneg64_69 in64_69 sn64_69 78000.000000
Rwneg64_70 in64_70 sn64_70 202000.000000
Rwneg64_71 in64_71 sn64_71 78000.000000
Rwneg64_72 in64_72 sn64_72 202000.000000
Rwneg64_73 in64_73 sn64_73 202000.000000
Rwneg64_74 in64_74 sn64_74 202000.000000
Rwneg64_75 in64_75 sn64_75 202000.000000
Rwneg64_76 in64_76 sn64_76 202000.000000
Rwneg64_77 in64_77 sn64_77 78000.000000
Rwneg64_78 in64_78 sn64_78 202000.000000
Rwneg64_79 in64_79 sn64_79 78000.000000
Rwneg64_80 in64_80 sn64_80 78000.000000
Rwneg64_81 in64_81 sn64_81 202000.000000
Rwneg64_82 in64_82 sn64_82 78000.000000
Rwneg64_83 in64_83 sn64_83 202000.000000
Rwneg64_84 in64_84 sn64_84 202000.000000
Rwneg65_1 in65_1 sn65_1 202000.000000
Rwneg65_2 in65_2 sn65_2 78000.000000
Rwneg65_3 in65_3 sn65_3 202000.000000
Rwneg65_4 in65_4 sn65_4 202000.000000
Rwneg65_5 in65_5 sn65_5 202000.000000
Rwneg65_6 in65_6 sn65_6 78000.000000
Rwneg65_7 in65_7 sn65_7 78000.000000
Rwneg65_8 in65_8 sn65_8 202000.000000
Rwneg65_9 in65_9 sn65_9 78000.000000
Rwneg65_10 in65_10 sn65_10 78000.000000
Rwneg65_11 in65_11 sn65_11 78000.000000
Rwneg65_12 in65_12 sn65_12 78000.000000
Rwneg65_13 in65_13 sn65_13 202000.000000
Rwneg65_14 in65_14 sn65_14 202000.000000
Rwneg65_15 in65_15 sn65_15 78000.000000
Rwneg65_16 in65_16 sn65_16 78000.000000
Rwneg65_17 in65_17 sn65_17 78000.000000
Rwneg65_18 in65_18 sn65_18 202000.000000
Rwneg65_19 in65_19 sn65_19 202000.000000
Rwneg65_20 in65_20 sn65_20 202000.000000
Rwneg65_21 in65_21 sn65_21 78000.000000
Rwneg65_22 in65_22 sn65_22 78000.000000
Rwneg65_23 in65_23 sn65_23 202000.000000
Rwneg65_24 in65_24 sn65_24 78000.000000
Rwneg65_25 in65_25 sn65_25 202000.000000
Rwneg65_26 in65_26 sn65_26 202000.000000
Rwneg65_27 in65_27 sn65_27 202000.000000
Rwneg65_28 in65_28 sn65_28 202000.000000
Rwneg65_29 in65_29 sn65_29 78000.000000
Rwneg65_30 in65_30 sn65_30 202000.000000
Rwneg65_31 in65_31 sn65_31 202000.000000
Rwneg65_32 in65_32 sn65_32 202000.000000
Rwneg65_33 in65_33 sn65_33 202000.000000
Rwneg65_34 in65_34 sn65_34 78000.000000
Rwneg65_35 in65_35 sn65_35 202000.000000
Rwneg65_36 in65_36 sn65_36 78000.000000
Rwneg65_37 in65_37 sn65_37 202000.000000
Rwneg65_38 in65_38 sn65_38 202000.000000
Rwneg65_39 in65_39 sn65_39 78000.000000
Rwneg65_40 in65_40 sn65_40 202000.000000
Rwneg65_41 in65_41 sn65_41 78000.000000
Rwneg65_42 in65_42 sn65_42 202000.000000
Rwneg65_43 in65_43 sn65_43 202000.000000
Rwneg65_44 in65_44 sn65_44 78000.000000
Rwneg65_45 in65_45 sn65_45 202000.000000
Rwneg65_46 in65_46 sn65_46 202000.000000
Rwneg65_47 in65_47 sn65_47 78000.000000
Rwneg65_48 in65_48 sn65_48 78000.000000
Rwneg65_49 in65_49 sn65_49 202000.000000
Rwneg65_50 in65_50 sn65_50 202000.000000
Rwneg65_51 in65_51 sn65_51 202000.000000
Rwneg65_52 in65_52 sn65_52 202000.000000
Rwneg65_53 in65_53 sn65_53 202000.000000
Rwneg65_54 in65_54 sn65_54 202000.000000
Rwneg65_55 in65_55 sn65_55 78000.000000
Rwneg65_56 in65_56 sn65_56 202000.000000
Rwneg65_57 in65_57 sn65_57 78000.000000
Rwneg65_58 in65_58 sn65_58 78000.000000
Rwneg65_59 in65_59 sn65_59 202000.000000
Rwneg65_60 in65_60 sn65_60 78000.000000
Rwneg65_61 in65_61 sn65_61 78000.000000
Rwneg65_62 in65_62 sn65_62 202000.000000
Rwneg65_63 in65_63 sn65_63 78000.000000
Rwneg65_64 in65_64 sn65_64 78000.000000
Rwneg65_65 in65_65 sn65_65 78000.000000
Rwneg65_66 in65_66 sn65_66 202000.000000
Rwneg65_67 in65_67 sn65_67 202000.000000
Rwneg65_68 in65_68 sn65_68 78000.000000
Rwneg65_69 in65_69 sn65_69 78000.000000
Rwneg65_70 in65_70 sn65_70 78000.000000
Rwneg65_71 in65_71 sn65_71 78000.000000
Rwneg65_72 in65_72 sn65_72 78000.000000
Rwneg65_73 in65_73 sn65_73 78000.000000
Rwneg65_74 in65_74 sn65_74 202000.000000
Rwneg65_75 in65_75 sn65_75 202000.000000
Rwneg65_76 in65_76 sn65_76 78000.000000
Rwneg65_77 in65_77 sn65_77 202000.000000
Rwneg65_78 in65_78 sn65_78 202000.000000
Rwneg65_79 in65_79 sn65_79 78000.000000
Rwneg65_80 in65_80 sn65_80 202000.000000
Rwneg65_81 in65_81 sn65_81 78000.000000
Rwneg65_82 in65_82 sn65_82 78000.000000
Rwneg65_83 in65_83 sn65_83 202000.000000
Rwneg65_84 in65_84 sn65_84 202000.000000
Rwneg66_1 in66_1 sn66_1 202000.000000
Rwneg66_2 in66_2 sn66_2 78000.000000
Rwneg66_3 in66_3 sn66_3 202000.000000
Rwneg66_4 in66_4 sn66_4 78000.000000
Rwneg66_5 in66_5 sn66_5 202000.000000
Rwneg66_6 in66_6 sn66_6 78000.000000
Rwneg66_7 in66_7 sn66_7 202000.000000
Rwneg66_8 in66_8 sn66_8 78000.000000
Rwneg66_9 in66_9 sn66_9 202000.000000
Rwneg66_10 in66_10 sn66_10 78000.000000
Rwneg66_11 in66_11 sn66_11 78000.000000
Rwneg66_12 in66_12 sn66_12 78000.000000
Rwneg66_13 in66_13 sn66_13 78000.000000
Rwneg66_14 in66_14 sn66_14 202000.000000
Rwneg66_15 in66_15 sn66_15 202000.000000
Rwneg66_16 in66_16 sn66_16 202000.000000
Rwneg66_17 in66_17 sn66_17 78000.000000
Rwneg66_18 in66_18 sn66_18 78000.000000
Rwneg66_19 in66_19 sn66_19 78000.000000
Rwneg66_20 in66_20 sn66_20 202000.000000
Rwneg66_21 in66_21 sn66_21 202000.000000
Rwneg66_22 in66_22 sn66_22 78000.000000
Rwneg66_23 in66_23 sn66_23 78000.000000
Rwneg66_24 in66_24 sn66_24 202000.000000
Rwneg66_25 in66_25 sn66_25 78000.000000
Rwneg66_26 in66_26 sn66_26 202000.000000
Rwneg66_27 in66_27 sn66_27 78000.000000
Rwneg66_28 in66_28 sn66_28 202000.000000
Rwneg66_29 in66_29 sn66_29 202000.000000
Rwneg66_30 in66_30 sn66_30 202000.000000
Rwneg66_31 in66_31 sn66_31 78000.000000
Rwneg66_32 in66_32 sn66_32 78000.000000
Rwneg66_33 in66_33 sn66_33 202000.000000
Rwneg66_34 in66_34 sn66_34 78000.000000
Rwneg66_35 in66_35 sn66_35 202000.000000
Rwneg66_36 in66_36 sn66_36 78000.000000
Rwneg66_37 in66_37 sn66_37 202000.000000
Rwneg66_38 in66_38 sn66_38 78000.000000
Rwneg66_39 in66_39 sn66_39 78000.000000
Rwneg66_40 in66_40 sn66_40 78000.000000
Rwneg66_41 in66_41 sn66_41 202000.000000
Rwneg66_42 in66_42 sn66_42 202000.000000
Rwneg66_43 in66_43 sn66_43 202000.000000
Rwneg66_44 in66_44 sn66_44 202000.000000
Rwneg66_45 in66_45 sn66_45 78000.000000
Rwneg66_46 in66_46 sn66_46 78000.000000
Rwneg66_47 in66_47 sn66_47 78000.000000
Rwneg66_48 in66_48 sn66_48 78000.000000
Rwneg66_49 in66_49 sn66_49 202000.000000
Rwneg66_50 in66_50 sn66_50 202000.000000
Rwneg66_51 in66_51 sn66_51 202000.000000
Rwneg66_52 in66_52 sn66_52 202000.000000
Rwneg66_53 in66_53 sn66_53 78000.000000
Rwneg66_54 in66_54 sn66_54 202000.000000
Rwneg66_55 in66_55 sn66_55 202000.000000
Rwneg66_56 in66_56 sn66_56 78000.000000
Rwneg66_57 in66_57 sn66_57 202000.000000
Rwneg66_58 in66_58 sn66_58 78000.000000
Rwneg66_59 in66_59 sn66_59 202000.000000
Rwneg66_60 in66_60 sn66_60 78000.000000
Rwneg66_61 in66_61 sn66_61 202000.000000
Rwneg66_62 in66_62 sn66_62 202000.000000
Rwneg66_63 in66_63 sn66_63 202000.000000
Rwneg66_64 in66_64 sn66_64 78000.000000
Rwneg66_65 in66_65 sn66_65 202000.000000
Rwneg66_66 in66_66 sn66_66 202000.000000
Rwneg66_67 in66_67 sn66_67 78000.000000
Rwneg66_68 in66_68 sn66_68 78000.000000
Rwneg66_69 in66_69 sn66_69 78000.000000
Rwneg66_70 in66_70 sn66_70 202000.000000
Rwneg66_71 in66_71 sn66_71 78000.000000
Rwneg66_72 in66_72 sn66_72 202000.000000
Rwneg66_73 in66_73 sn66_73 78000.000000
Rwneg66_74 in66_74 sn66_74 78000.000000
Rwneg66_75 in66_75 sn66_75 78000.000000
Rwneg66_76 in66_76 sn66_76 202000.000000
Rwneg66_77 in66_77 sn66_77 78000.000000
Rwneg66_78 in66_78 sn66_78 78000.000000
Rwneg66_79 in66_79 sn66_79 78000.000000
Rwneg66_80 in66_80 sn66_80 202000.000000
Rwneg66_81 in66_81 sn66_81 202000.000000
Rwneg66_82 in66_82 sn66_82 202000.000000
Rwneg66_83 in66_83 sn66_83 78000.000000
Rwneg66_84 in66_84 sn66_84 202000.000000
Rwneg67_1 in67_1 sn67_1 78000.000000
Rwneg67_2 in67_2 sn67_2 78000.000000
Rwneg67_3 in67_3 sn67_3 202000.000000
Rwneg67_4 in67_4 sn67_4 78000.000000
Rwneg67_5 in67_5 sn67_5 202000.000000
Rwneg67_6 in67_6 sn67_6 78000.000000
Rwneg67_7 in67_7 sn67_7 202000.000000
Rwneg67_8 in67_8 sn67_8 78000.000000
Rwneg67_9 in67_9 sn67_9 78000.000000
Rwneg67_10 in67_10 sn67_10 202000.000000
Rwneg67_11 in67_11 sn67_11 78000.000000
Rwneg67_12 in67_12 sn67_12 78000.000000
Rwneg67_13 in67_13 sn67_13 78000.000000
Rwneg67_14 in67_14 sn67_14 78000.000000
Rwneg67_15 in67_15 sn67_15 78000.000000
Rwneg67_16 in67_16 sn67_16 202000.000000
Rwneg67_17 in67_17 sn67_17 202000.000000
Rwneg67_18 in67_18 sn67_18 78000.000000
Rwneg67_19 in67_19 sn67_19 202000.000000
Rwneg67_20 in67_20 sn67_20 78000.000000
Rwneg67_21 in67_21 sn67_21 202000.000000
Rwneg67_22 in67_22 sn67_22 202000.000000
Rwneg67_23 in67_23 sn67_23 202000.000000
Rwneg67_24 in67_24 sn67_24 202000.000000
Rwneg67_25 in67_25 sn67_25 78000.000000
Rwneg67_26 in67_26 sn67_26 78000.000000
Rwneg67_27 in67_27 sn67_27 202000.000000
Rwneg67_28 in67_28 sn67_28 202000.000000
Rwneg67_29 in67_29 sn67_29 202000.000000
Rwneg67_30 in67_30 sn67_30 202000.000000
Rwneg67_31 in67_31 sn67_31 202000.000000
Rwneg67_32 in67_32 sn67_32 202000.000000
Rwneg67_33 in67_33 sn67_33 202000.000000
Rwneg67_34 in67_34 sn67_34 78000.000000
Rwneg67_35 in67_35 sn67_35 78000.000000
Rwneg67_36 in67_36 sn67_36 78000.000000
Rwneg67_37 in67_37 sn67_37 202000.000000
Rwneg67_38 in67_38 sn67_38 202000.000000
Rwneg67_39 in67_39 sn67_39 78000.000000
Rwneg67_40 in67_40 sn67_40 78000.000000
Rwneg67_41 in67_41 sn67_41 78000.000000
Rwneg67_42 in67_42 sn67_42 78000.000000
Rwneg67_43 in67_43 sn67_43 78000.000000
Rwneg67_44 in67_44 sn67_44 202000.000000
Rwneg67_45 in67_45 sn67_45 202000.000000
Rwneg67_46 in67_46 sn67_46 202000.000000
Rwneg67_47 in67_47 sn67_47 78000.000000
Rwneg67_48 in67_48 sn67_48 202000.000000
Rwneg67_49 in67_49 sn67_49 78000.000000
Rwneg67_50 in67_50 sn67_50 78000.000000
Rwneg67_51 in67_51 sn67_51 202000.000000
Rwneg67_52 in67_52 sn67_52 78000.000000
Rwneg67_53 in67_53 sn67_53 78000.000000
Rwneg67_54 in67_54 sn67_54 202000.000000
Rwneg67_55 in67_55 sn67_55 202000.000000
Rwneg67_56 in67_56 sn67_56 78000.000000
Rwneg67_57 in67_57 sn67_57 202000.000000
Rwneg67_58 in67_58 sn67_58 202000.000000
Rwneg67_59 in67_59 sn67_59 202000.000000
Rwneg67_60 in67_60 sn67_60 78000.000000
Rwneg67_61 in67_61 sn67_61 202000.000000
Rwneg67_62 in67_62 sn67_62 202000.000000
Rwneg67_63 in67_63 sn67_63 78000.000000
Rwneg67_64 in67_64 sn67_64 202000.000000
Rwneg67_65 in67_65 sn67_65 78000.000000
Rwneg67_66 in67_66 sn67_66 78000.000000
Rwneg67_67 in67_67 sn67_67 202000.000000
Rwneg67_68 in67_68 sn67_68 78000.000000
Rwneg67_69 in67_69 sn67_69 78000.000000
Rwneg67_70 in67_70 sn67_70 202000.000000
Rwneg67_71 in67_71 sn67_71 78000.000000
Rwneg67_72 in67_72 sn67_72 202000.000000
Rwneg67_73 in67_73 sn67_73 202000.000000
Rwneg67_74 in67_74 sn67_74 202000.000000
Rwneg67_75 in67_75 sn67_75 202000.000000
Rwneg67_76 in67_76 sn67_76 78000.000000
Rwneg67_77 in67_77 sn67_77 202000.000000
Rwneg67_78 in67_78 sn67_78 202000.000000
Rwneg67_79 in67_79 sn67_79 78000.000000
Rwneg67_80 in67_80 sn67_80 202000.000000
Rwneg67_81 in67_81 sn67_81 202000.000000
Rwneg67_82 in67_82 sn67_82 78000.000000
Rwneg67_83 in67_83 sn67_83 202000.000000
Rwneg67_84 in67_84 sn67_84 78000.000000
Rwneg68_1 in68_1 sn68_1 202000.000000
Rwneg68_2 in68_2 sn68_2 202000.000000
Rwneg68_3 in68_3 sn68_3 202000.000000
Rwneg68_4 in68_4 sn68_4 78000.000000
Rwneg68_5 in68_5 sn68_5 78000.000000
Rwneg68_6 in68_6 sn68_6 202000.000000
Rwneg68_7 in68_7 sn68_7 78000.000000
Rwneg68_8 in68_8 sn68_8 78000.000000
Rwneg68_9 in68_9 sn68_9 78000.000000
Rwneg68_10 in68_10 sn68_10 202000.000000
Rwneg68_11 in68_11 sn68_11 78000.000000
Rwneg68_12 in68_12 sn68_12 78000.000000
Rwneg68_13 in68_13 sn68_13 78000.000000
Rwneg68_14 in68_14 sn68_14 202000.000000
Rwneg68_15 in68_15 sn68_15 78000.000000
Rwneg68_16 in68_16 sn68_16 78000.000000
Rwneg68_17 in68_17 sn68_17 78000.000000
Rwneg68_18 in68_18 sn68_18 202000.000000
Rwneg68_19 in68_19 sn68_19 202000.000000
Rwneg68_20 in68_20 sn68_20 202000.000000
Rwneg68_21 in68_21 sn68_21 202000.000000
Rwneg68_22 in68_22 sn68_22 202000.000000
Rwneg68_23 in68_23 sn68_23 78000.000000
Rwneg68_24 in68_24 sn68_24 202000.000000
Rwneg68_25 in68_25 sn68_25 78000.000000
Rwneg68_26 in68_26 sn68_26 202000.000000
Rwneg68_27 in68_27 sn68_27 202000.000000
Rwneg68_28 in68_28 sn68_28 202000.000000
Rwneg68_29 in68_29 sn68_29 78000.000000
Rwneg68_30 in68_30 sn68_30 78000.000000
Rwneg68_31 in68_31 sn68_31 78000.000000
Rwneg68_32 in68_32 sn68_32 202000.000000
Rwneg68_33 in68_33 sn68_33 202000.000000
Rwneg68_34 in68_34 sn68_34 78000.000000
Rwneg68_35 in68_35 sn68_35 202000.000000
Rwneg68_36 in68_36 sn68_36 202000.000000
Rwneg68_37 in68_37 sn68_37 202000.000000
Rwneg68_38 in68_38 sn68_38 202000.000000
Rwneg68_39 in68_39 sn68_39 78000.000000
Rwneg68_40 in68_40 sn68_40 78000.000000
Rwneg68_41 in68_41 sn68_41 78000.000000
Rwneg68_42 in68_42 sn68_42 202000.000000
Rwneg68_43 in68_43 sn68_43 202000.000000
Rwneg68_44 in68_44 sn68_44 202000.000000
Rwneg68_45 in68_45 sn68_45 202000.000000
Rwneg68_46 in68_46 sn68_46 78000.000000
Rwneg68_47 in68_47 sn68_47 78000.000000
Rwneg68_48 in68_48 sn68_48 78000.000000
Rwneg68_49 in68_49 sn68_49 78000.000000
Rwneg68_50 in68_50 sn68_50 202000.000000
Rwneg68_51 in68_51 sn68_51 202000.000000
Rwneg68_52 in68_52 sn68_52 202000.000000
Rwneg68_53 in68_53 sn68_53 78000.000000
Rwneg68_54 in68_54 sn68_54 78000.000000
Rwneg68_55 in68_55 sn68_55 78000.000000
Rwneg68_56 in68_56 sn68_56 78000.000000
Rwneg68_57 in68_57 sn68_57 202000.000000
Rwneg68_58 in68_58 sn68_58 78000.000000
Rwneg68_59 in68_59 sn68_59 202000.000000
Rwneg68_60 in68_60 sn68_60 78000.000000
Rwneg68_61 in68_61 sn68_61 202000.000000
Rwneg68_62 in68_62 sn68_62 78000.000000
Rwneg68_63 in68_63 sn68_63 78000.000000
Rwneg68_64 in68_64 sn68_64 202000.000000
Rwneg68_65 in68_65 sn68_65 78000.000000
Rwneg68_66 in68_66 sn68_66 78000.000000
Rwneg68_67 in68_67 sn68_67 202000.000000
Rwneg68_68 in68_68 sn68_68 78000.000000
Rwneg68_69 in68_69 sn68_69 78000.000000
Rwneg68_70 in68_70 sn68_70 78000.000000
Rwneg68_71 in68_71 sn68_71 78000.000000
Rwneg68_72 in68_72 sn68_72 202000.000000
Rwneg68_73 in68_73 sn68_73 78000.000000
Rwneg68_74 in68_74 sn68_74 78000.000000
Rwneg68_75 in68_75 sn68_75 202000.000000
Rwneg68_76 in68_76 sn68_76 78000.000000
Rwneg68_77 in68_77 sn68_77 202000.000000
Rwneg68_78 in68_78 sn68_78 202000.000000
Rwneg68_79 in68_79 sn68_79 78000.000000
Rwneg68_80 in68_80 sn68_80 78000.000000
Rwneg68_81 in68_81 sn68_81 78000.000000
Rwneg68_82 in68_82 sn68_82 78000.000000
Rwneg68_83 in68_83 sn68_83 202000.000000
Rwneg68_84 in68_84 sn68_84 202000.000000
Rwneg69_1 in69_1 sn69_1 202000.000000
Rwneg69_2 in69_2 sn69_2 78000.000000
Rwneg69_3 in69_3 sn69_3 78000.000000
Rwneg69_4 in69_4 sn69_4 202000.000000
Rwneg69_5 in69_5 sn69_5 202000.000000
Rwneg69_6 in69_6 sn69_6 202000.000000
Rwneg69_7 in69_7 sn69_7 78000.000000
Rwneg69_8 in69_8 sn69_8 78000.000000
Rwneg69_9 in69_9 sn69_9 202000.000000
Rwneg69_10 in69_10 sn69_10 202000.000000
Rwneg69_11 in69_11 sn69_11 78000.000000
Rwneg69_12 in69_12 sn69_12 202000.000000
Rwneg69_13 in69_13 sn69_13 202000.000000
Rwneg69_14 in69_14 sn69_14 78000.000000
Rwneg69_15 in69_15 sn69_15 78000.000000
Rwneg69_16 in69_16 sn69_16 202000.000000
Rwneg69_17 in69_17 sn69_17 78000.000000
Rwneg69_18 in69_18 sn69_18 202000.000000
Rwneg69_19 in69_19 sn69_19 202000.000000
Rwneg69_20 in69_20 sn69_20 202000.000000
Rwneg69_21 in69_21 sn69_21 78000.000000
Rwneg69_22 in69_22 sn69_22 78000.000000
Rwneg69_23 in69_23 sn69_23 202000.000000
Rwneg69_24 in69_24 sn69_24 202000.000000
Rwneg69_25 in69_25 sn69_25 78000.000000
Rwneg69_26 in69_26 sn69_26 78000.000000
Rwneg69_27 in69_27 sn69_27 202000.000000
Rwneg69_28 in69_28 sn69_28 202000.000000
Rwneg69_29 in69_29 sn69_29 78000.000000
Rwneg69_30 in69_30 sn69_30 78000.000000
Rwneg69_31 in69_31 sn69_31 78000.000000
Rwneg69_32 in69_32 sn69_32 202000.000000
Rwneg69_33 in69_33 sn69_33 78000.000000
Rwneg69_34 in69_34 sn69_34 202000.000000
Rwneg69_35 in69_35 sn69_35 78000.000000
Rwneg69_36 in69_36 sn69_36 202000.000000
Rwneg69_37 in69_37 sn69_37 78000.000000
Rwneg69_38 in69_38 sn69_38 202000.000000
Rwneg69_39 in69_39 sn69_39 202000.000000
Rwneg69_40 in69_40 sn69_40 202000.000000
Rwneg69_41 in69_41 sn69_41 78000.000000
Rwneg69_42 in69_42 sn69_42 78000.000000
Rwneg69_43 in69_43 sn69_43 202000.000000
Rwneg69_44 in69_44 sn69_44 78000.000000
Rwneg69_45 in69_45 sn69_45 202000.000000
Rwneg69_46 in69_46 sn69_46 78000.000000
Rwneg69_47 in69_47 sn69_47 202000.000000
Rwneg69_48 in69_48 sn69_48 202000.000000
Rwneg69_49 in69_49 sn69_49 78000.000000
Rwneg69_50 in69_50 sn69_50 78000.000000
Rwneg69_51 in69_51 sn69_51 78000.000000
Rwneg69_52 in69_52 sn69_52 78000.000000
Rwneg69_53 in69_53 sn69_53 78000.000000
Rwneg69_54 in69_54 sn69_54 202000.000000
Rwneg69_55 in69_55 sn69_55 78000.000000
Rwneg69_56 in69_56 sn69_56 202000.000000
Rwneg69_57 in69_57 sn69_57 202000.000000
Rwneg69_58 in69_58 sn69_58 78000.000000
Rwneg69_59 in69_59 sn69_59 78000.000000
Rwneg69_60 in69_60 sn69_60 78000.000000
Rwneg69_61 in69_61 sn69_61 78000.000000
Rwneg69_62 in69_62 sn69_62 78000.000000
Rwneg69_63 in69_63 sn69_63 202000.000000
Rwneg69_64 in69_64 sn69_64 78000.000000
Rwneg69_65 in69_65 sn69_65 202000.000000
Rwneg69_66 in69_66 sn69_66 202000.000000
Rwneg69_67 in69_67 sn69_67 202000.000000
Rwneg69_68 in69_68 sn69_68 202000.000000
Rwneg69_69 in69_69 sn69_69 202000.000000
Rwneg69_70 in69_70 sn69_70 202000.000000
Rwneg69_71 in69_71 sn69_71 202000.000000
Rwneg69_72 in69_72 sn69_72 78000.000000
Rwneg69_73 in69_73 sn69_73 202000.000000
Rwneg69_74 in69_74 sn69_74 78000.000000
Rwneg69_75 in69_75 sn69_75 202000.000000
Rwneg69_76 in69_76 sn69_76 202000.000000
Rwneg69_77 in69_77 sn69_77 202000.000000
Rwneg69_78 in69_78 sn69_78 78000.000000
Rwneg69_79 in69_79 sn69_79 202000.000000
Rwneg69_80 in69_80 sn69_80 202000.000000
Rwneg69_81 in69_81 sn69_81 202000.000000
Rwneg69_82 in69_82 sn69_82 202000.000000
Rwneg69_83 in69_83 sn69_83 78000.000000
Rwneg69_84 in69_84 sn69_84 202000.000000
Rwneg70_1 in70_1 sn70_1 202000.000000
Rwneg70_2 in70_2 sn70_2 202000.000000
Rwneg70_3 in70_3 sn70_3 78000.000000
Rwneg70_4 in70_4 sn70_4 78000.000000
Rwneg70_5 in70_5 sn70_5 202000.000000
Rwneg70_6 in70_6 sn70_6 202000.000000
Rwneg70_7 in70_7 sn70_7 202000.000000
Rwneg70_8 in70_8 sn70_8 202000.000000
Rwneg70_9 in70_9 sn70_9 202000.000000
Rwneg70_10 in70_10 sn70_10 78000.000000
Rwneg70_11 in70_11 sn70_11 78000.000000
Rwneg70_12 in70_12 sn70_12 202000.000000
Rwneg70_13 in70_13 sn70_13 78000.000000
Rwneg70_14 in70_14 sn70_14 202000.000000
Rwneg70_15 in70_15 sn70_15 202000.000000
Rwneg70_16 in70_16 sn70_16 78000.000000
Rwneg70_17 in70_17 sn70_17 78000.000000
Rwneg70_18 in70_18 sn70_18 202000.000000
Rwneg70_19 in70_19 sn70_19 202000.000000
Rwneg70_20 in70_20 sn70_20 202000.000000
Rwneg70_21 in70_21 sn70_21 78000.000000
Rwneg70_22 in70_22 sn70_22 78000.000000
Rwneg70_23 in70_23 sn70_23 202000.000000
Rwneg70_24 in70_24 sn70_24 78000.000000
Rwneg70_25 in70_25 sn70_25 202000.000000
Rwneg70_26 in70_26 sn70_26 202000.000000
Rwneg70_27 in70_27 sn70_27 202000.000000
Rwneg70_28 in70_28 sn70_28 78000.000000
Rwneg70_29 in70_29 sn70_29 202000.000000
Rwneg70_30 in70_30 sn70_30 78000.000000
Rwneg70_31 in70_31 sn70_31 78000.000000
Rwneg70_32 in70_32 sn70_32 78000.000000
Rwneg70_33 in70_33 sn70_33 78000.000000
Rwneg70_34 in70_34 sn70_34 202000.000000
Rwneg70_35 in70_35 sn70_35 78000.000000
Rwneg70_36 in70_36 sn70_36 78000.000000
Rwneg70_37 in70_37 sn70_37 202000.000000
Rwneg70_38 in70_38 sn70_38 78000.000000
Rwneg70_39 in70_39 sn70_39 202000.000000
Rwneg70_40 in70_40 sn70_40 202000.000000
Rwneg70_41 in70_41 sn70_41 78000.000000
Rwneg70_42 in70_42 sn70_42 202000.000000
Rwneg70_43 in70_43 sn70_43 202000.000000
Rwneg70_44 in70_44 sn70_44 78000.000000
Rwneg70_45 in70_45 sn70_45 202000.000000
Rwneg70_46 in70_46 sn70_46 202000.000000
Rwneg70_47 in70_47 sn70_47 78000.000000
Rwneg70_48 in70_48 sn70_48 202000.000000
Rwneg70_49 in70_49 sn70_49 202000.000000
Rwneg70_50 in70_50 sn70_50 202000.000000
Rwneg70_51 in70_51 sn70_51 78000.000000
Rwneg70_52 in70_52 sn70_52 202000.000000
Rwneg70_53 in70_53 sn70_53 202000.000000
Rwneg70_54 in70_54 sn70_54 202000.000000
Rwneg70_55 in70_55 sn70_55 78000.000000
Rwneg70_56 in70_56 sn70_56 202000.000000
Rwneg70_57 in70_57 sn70_57 78000.000000
Rwneg70_58 in70_58 sn70_58 202000.000000
Rwneg70_59 in70_59 sn70_59 78000.000000
Rwneg70_60 in70_60 sn70_60 202000.000000
Rwneg70_61 in70_61 sn70_61 78000.000000
Rwneg70_62 in70_62 sn70_62 78000.000000
Rwneg70_63 in70_63 sn70_63 202000.000000
Rwneg70_64 in70_64 sn70_64 202000.000000
Rwneg70_65 in70_65 sn70_65 202000.000000
Rwneg70_66 in70_66 sn70_66 202000.000000
Rwneg70_67 in70_67 sn70_67 202000.000000
Rwneg70_68 in70_68 sn70_68 78000.000000
Rwneg70_69 in70_69 sn70_69 202000.000000
Rwneg70_70 in70_70 sn70_70 78000.000000
Rwneg70_71 in70_71 sn70_71 202000.000000
Rwneg70_72 in70_72 sn70_72 202000.000000
Rwneg70_73 in70_73 sn70_73 202000.000000
Rwneg70_74 in70_74 sn70_74 202000.000000
Rwneg70_75 in70_75 sn70_75 78000.000000
Rwneg70_76 in70_76 sn70_76 202000.000000
Rwneg70_77 in70_77 sn70_77 78000.000000
Rwneg70_78 in70_78 sn70_78 202000.000000
Rwneg70_79 in70_79 sn70_79 202000.000000
Rwneg70_80 in70_80 sn70_80 202000.000000
Rwneg70_81 in70_81 sn70_81 78000.000000
Rwneg70_82 in70_82 sn70_82 202000.000000
Rwneg70_83 in70_83 sn70_83 202000.000000
Rwneg70_84 in70_84 sn70_84 78000.000000
Rwneg71_1 in71_1 sn71_1 202000.000000
Rwneg71_2 in71_2 sn71_2 78000.000000
Rwneg71_3 in71_3 sn71_3 202000.000000
Rwneg71_4 in71_4 sn71_4 202000.000000
Rwneg71_5 in71_5 sn71_5 78000.000000
Rwneg71_6 in71_6 sn71_6 202000.000000
Rwneg71_7 in71_7 sn71_7 78000.000000
Rwneg71_8 in71_8 sn71_8 78000.000000
Rwneg71_9 in71_9 sn71_9 202000.000000
Rwneg71_10 in71_10 sn71_10 78000.000000
Rwneg71_11 in71_11 sn71_11 78000.000000
Rwneg71_12 in71_12 sn71_12 202000.000000
Rwneg71_13 in71_13 sn71_13 78000.000000
Rwneg71_14 in71_14 sn71_14 202000.000000
Rwneg71_15 in71_15 sn71_15 202000.000000
Rwneg71_16 in71_16 sn71_16 202000.000000
Rwneg71_17 in71_17 sn71_17 202000.000000
Rwneg71_18 in71_18 sn71_18 78000.000000
Rwneg71_19 in71_19 sn71_19 202000.000000
Rwneg71_20 in71_20 sn71_20 78000.000000
Rwneg71_21 in71_21 sn71_21 78000.000000
Rwneg71_22 in71_22 sn71_22 202000.000000
Rwneg71_23 in71_23 sn71_23 78000.000000
Rwneg71_24 in71_24 sn71_24 202000.000000
Rwneg71_25 in71_25 sn71_25 202000.000000
Rwneg71_26 in71_26 sn71_26 202000.000000
Rwneg71_27 in71_27 sn71_27 78000.000000
Rwneg71_28 in71_28 sn71_28 78000.000000
Rwneg71_29 in71_29 sn71_29 78000.000000
Rwneg71_30 in71_30 sn71_30 202000.000000
Rwneg71_31 in71_31 sn71_31 202000.000000
Rwneg71_32 in71_32 sn71_32 202000.000000
Rwneg71_33 in71_33 sn71_33 78000.000000
Rwneg71_34 in71_34 sn71_34 202000.000000
Rwneg71_35 in71_35 sn71_35 202000.000000
Rwneg71_36 in71_36 sn71_36 202000.000000
Rwneg71_37 in71_37 sn71_37 78000.000000
Rwneg71_38 in71_38 sn71_38 202000.000000
Rwneg71_39 in71_39 sn71_39 202000.000000
Rwneg71_40 in71_40 sn71_40 202000.000000
Rwneg71_41 in71_41 sn71_41 202000.000000
Rwneg71_42 in71_42 sn71_42 78000.000000
Rwneg71_43 in71_43 sn71_43 78000.000000
Rwneg71_44 in71_44 sn71_44 202000.000000
Rwneg71_45 in71_45 sn71_45 78000.000000
Rwneg71_46 in71_46 sn71_46 202000.000000
Rwneg71_47 in71_47 sn71_47 202000.000000
Rwneg71_48 in71_48 sn71_48 202000.000000
Rwneg71_49 in71_49 sn71_49 202000.000000
Rwneg71_50 in71_50 sn71_50 202000.000000
Rwneg71_51 in71_51 sn71_51 202000.000000
Rwneg71_52 in71_52 sn71_52 202000.000000
Rwneg71_53 in71_53 sn71_53 78000.000000
Rwneg71_54 in71_54 sn71_54 78000.000000
Rwneg71_55 in71_55 sn71_55 78000.000000
Rwneg71_56 in71_56 sn71_56 78000.000000
Rwneg71_57 in71_57 sn71_57 202000.000000
Rwneg71_58 in71_58 sn71_58 202000.000000
Rwneg71_59 in71_59 sn71_59 78000.000000
Rwneg71_60 in71_60 sn71_60 202000.000000
Rwneg71_61 in71_61 sn71_61 202000.000000
Rwneg71_62 in71_62 sn71_62 78000.000000
Rwneg71_63 in71_63 sn71_63 202000.000000
Rwneg71_64 in71_64 sn71_64 78000.000000
Rwneg71_65 in71_65 sn71_65 78000.000000
Rwneg71_66 in71_66 sn71_66 202000.000000
Rwneg71_67 in71_67 sn71_67 202000.000000
Rwneg71_68 in71_68 sn71_68 202000.000000
Rwneg71_69 in71_69 sn71_69 78000.000000
Rwneg71_70 in71_70 sn71_70 202000.000000
Rwneg71_71 in71_71 sn71_71 202000.000000
Rwneg71_72 in71_72 sn71_72 202000.000000
Rwneg71_73 in71_73 sn71_73 202000.000000
Rwneg71_74 in71_74 sn71_74 202000.000000
Rwneg71_75 in71_75 sn71_75 202000.000000
Rwneg71_76 in71_76 sn71_76 202000.000000
Rwneg71_77 in71_77 sn71_77 202000.000000
Rwneg71_78 in71_78 sn71_78 78000.000000
Rwneg71_79 in71_79 sn71_79 78000.000000
Rwneg71_80 in71_80 sn71_80 78000.000000
Rwneg71_81 in71_81 sn71_81 78000.000000
Rwneg71_82 in71_82 sn71_82 78000.000000
Rwneg71_83 in71_83 sn71_83 202000.000000
Rwneg71_84 in71_84 sn71_84 202000.000000
Rwneg72_1 in72_1 sn72_1 202000.000000
Rwneg72_2 in72_2 sn72_2 78000.000000
Rwneg72_3 in72_3 sn72_3 78000.000000
Rwneg72_4 in72_4 sn72_4 78000.000000
Rwneg72_5 in72_5 sn72_5 78000.000000
Rwneg72_6 in72_6 sn72_6 202000.000000
Rwneg72_7 in72_7 sn72_7 78000.000000
Rwneg72_8 in72_8 sn72_8 78000.000000
Rwneg72_9 in72_9 sn72_9 78000.000000
Rwneg72_10 in72_10 sn72_10 202000.000000
Rwneg72_11 in72_11 sn72_11 202000.000000
Rwneg72_12 in72_12 sn72_12 78000.000000
Rwneg72_13 in72_13 sn72_13 78000.000000
Rwneg72_14 in72_14 sn72_14 78000.000000
Rwneg72_15 in72_15 sn72_15 202000.000000
Rwneg72_16 in72_16 sn72_16 202000.000000
Rwneg72_17 in72_17 sn72_17 202000.000000
Rwneg72_18 in72_18 sn72_18 78000.000000
Rwneg72_19 in72_19 sn72_19 78000.000000
Rwneg72_20 in72_20 sn72_20 202000.000000
Rwneg72_21 in72_21 sn72_21 202000.000000
Rwneg72_22 in72_22 sn72_22 202000.000000
Rwneg72_23 in72_23 sn72_23 202000.000000
Rwneg72_24 in72_24 sn72_24 202000.000000
Rwneg72_25 in72_25 sn72_25 78000.000000
Rwneg72_26 in72_26 sn72_26 78000.000000
Rwneg72_27 in72_27 sn72_27 78000.000000
Rwneg72_28 in72_28 sn72_28 78000.000000
Rwneg72_29 in72_29 sn72_29 202000.000000
Rwneg72_30 in72_30 sn72_30 202000.000000
Rwneg72_31 in72_31 sn72_31 78000.000000
Rwneg72_32 in72_32 sn72_32 202000.000000
Rwneg72_33 in72_33 sn72_33 202000.000000
Rwneg72_34 in72_34 sn72_34 78000.000000
Rwneg72_35 in72_35 sn72_35 78000.000000
Rwneg72_36 in72_36 sn72_36 78000.000000
Rwneg72_37 in72_37 sn72_37 202000.000000
Rwneg72_38 in72_38 sn72_38 78000.000000
Rwneg72_39 in72_39 sn72_39 78000.000000
Rwneg72_40 in72_40 sn72_40 202000.000000
Rwneg72_41 in72_41 sn72_41 202000.000000
Rwneg72_42 in72_42 sn72_42 202000.000000
Rwneg72_43 in72_43 sn72_43 78000.000000
Rwneg72_44 in72_44 sn72_44 202000.000000
Rwneg72_45 in72_45 sn72_45 202000.000000
Rwneg72_46 in72_46 sn72_46 78000.000000
Rwneg72_47 in72_47 sn72_47 78000.000000
Rwneg72_48 in72_48 sn72_48 202000.000000
Rwneg72_49 in72_49 sn72_49 78000.000000
Rwneg72_50 in72_50 sn72_50 202000.000000
Rwneg72_51 in72_51 sn72_51 202000.000000
Rwneg72_52 in72_52 sn72_52 78000.000000
Rwneg72_53 in72_53 sn72_53 78000.000000
Rwneg72_54 in72_54 sn72_54 78000.000000
Rwneg72_55 in72_55 sn72_55 78000.000000
Rwneg72_56 in72_56 sn72_56 78000.000000
Rwneg72_57 in72_57 sn72_57 202000.000000
Rwneg72_58 in72_58 sn72_58 202000.000000
Rwneg72_59 in72_59 sn72_59 202000.000000
Rwneg72_60 in72_60 sn72_60 78000.000000
Rwneg72_61 in72_61 sn72_61 202000.000000
Rwneg72_62 in72_62 sn72_62 202000.000000
Rwneg72_63 in72_63 sn72_63 78000.000000
Rwneg72_64 in72_64 sn72_64 202000.000000
Rwneg72_65 in72_65 sn72_65 78000.000000
Rwneg72_66 in72_66 sn72_66 78000.000000
Rwneg72_67 in72_67 sn72_67 78000.000000
Rwneg72_68 in72_68 sn72_68 202000.000000
Rwneg72_69 in72_69 sn72_69 78000.000000
Rwneg72_70 in72_70 sn72_70 202000.000000
Rwneg72_71 in72_71 sn72_71 78000.000000
Rwneg72_72 in72_72 sn72_72 78000.000000
Rwneg72_73 in72_73 sn72_73 202000.000000
Rwneg72_74 in72_74 sn72_74 202000.000000
Rwneg72_75 in72_75 sn72_75 78000.000000
Rwneg72_76 in72_76 sn72_76 78000.000000
Rwneg72_77 in72_77 sn72_77 202000.000000
Rwneg72_78 in72_78 sn72_78 202000.000000
Rwneg72_79 in72_79 sn72_79 202000.000000
Rwneg72_80 in72_80 sn72_80 202000.000000
Rwneg72_81 in72_81 sn72_81 202000.000000
Rwneg72_82 in72_82 sn72_82 78000.000000
Rwneg72_83 in72_83 sn72_83 78000.000000
Rwneg72_84 in72_84 sn72_84 202000.000000
Rwneg73_1 in73_1 sn73_1 202000.000000
Rwneg73_2 in73_2 sn73_2 202000.000000
Rwneg73_3 in73_3 sn73_3 202000.000000
Rwneg73_4 in73_4 sn73_4 202000.000000
Rwneg73_5 in73_5 sn73_5 78000.000000
Rwneg73_6 in73_6 sn73_6 78000.000000
Rwneg73_7 in73_7 sn73_7 78000.000000
Rwneg73_8 in73_8 sn73_8 202000.000000
Rwneg73_9 in73_9 sn73_9 78000.000000
Rwneg73_10 in73_10 sn73_10 202000.000000
Rwneg73_11 in73_11 sn73_11 78000.000000
Rwneg73_12 in73_12 sn73_12 78000.000000
Rwneg73_13 in73_13 sn73_13 78000.000000
Rwneg73_14 in73_14 sn73_14 202000.000000
Rwneg73_15 in73_15 sn73_15 78000.000000
Rwneg73_16 in73_16 sn73_16 78000.000000
Rwneg73_17 in73_17 sn73_17 78000.000000
Rwneg73_18 in73_18 sn73_18 202000.000000
Rwneg73_19 in73_19 sn73_19 78000.000000
Rwneg73_20 in73_20 sn73_20 202000.000000
Rwneg73_21 in73_21 sn73_21 78000.000000
Rwneg73_22 in73_22 sn73_22 202000.000000
Rwneg73_23 in73_23 sn73_23 78000.000000
Rwneg73_24 in73_24 sn73_24 202000.000000
Rwneg73_25 in73_25 sn73_25 202000.000000
Rwneg73_26 in73_26 sn73_26 78000.000000
Rwneg73_27 in73_27 sn73_27 202000.000000
Rwneg73_28 in73_28 sn73_28 78000.000000
Rwneg73_29 in73_29 sn73_29 78000.000000
Rwneg73_30 in73_30 sn73_30 202000.000000
Rwneg73_31 in73_31 sn73_31 78000.000000
Rwneg73_32 in73_32 sn73_32 202000.000000
Rwneg73_33 in73_33 sn73_33 202000.000000
Rwneg73_34 in73_34 sn73_34 202000.000000
Rwneg73_35 in73_35 sn73_35 202000.000000
Rwneg73_36 in73_36 sn73_36 202000.000000
Rwneg73_37 in73_37 sn73_37 78000.000000
Rwneg73_38 in73_38 sn73_38 78000.000000
Rwneg73_39 in73_39 sn73_39 78000.000000
Rwneg73_40 in73_40 sn73_40 78000.000000
Rwneg73_41 in73_41 sn73_41 78000.000000
Rwneg73_42 in73_42 sn73_42 78000.000000
Rwneg73_43 in73_43 sn73_43 202000.000000
Rwneg73_44 in73_44 sn73_44 78000.000000
Rwneg73_45 in73_45 sn73_45 78000.000000
Rwneg73_46 in73_46 sn73_46 202000.000000
Rwneg73_47 in73_47 sn73_47 78000.000000
Rwneg73_48 in73_48 sn73_48 78000.000000
Rwneg73_49 in73_49 sn73_49 202000.000000
Rwneg73_50 in73_50 sn73_50 78000.000000
Rwneg73_51 in73_51 sn73_51 78000.000000
Rwneg73_52 in73_52 sn73_52 202000.000000
Rwneg73_53 in73_53 sn73_53 78000.000000
Rwneg73_54 in73_54 sn73_54 78000.000000
Rwneg73_55 in73_55 sn73_55 78000.000000
Rwneg73_56 in73_56 sn73_56 202000.000000
Rwneg73_57 in73_57 sn73_57 202000.000000
Rwneg73_58 in73_58 sn73_58 202000.000000
Rwneg73_59 in73_59 sn73_59 78000.000000
Rwneg73_60 in73_60 sn73_60 202000.000000
Rwneg73_61 in73_61 sn73_61 202000.000000
Rwneg73_62 in73_62 sn73_62 78000.000000
Rwneg73_63 in73_63 sn73_63 78000.000000
Rwneg73_64 in73_64 sn73_64 78000.000000
Rwneg73_65 in73_65 sn73_65 78000.000000
Rwneg73_66 in73_66 sn73_66 202000.000000
Rwneg73_67 in73_67 sn73_67 202000.000000
Rwneg73_68 in73_68 sn73_68 78000.000000
Rwneg73_69 in73_69 sn73_69 202000.000000
Rwneg73_70 in73_70 sn73_70 78000.000000
Rwneg73_71 in73_71 sn73_71 202000.000000
Rwneg73_72 in73_72 sn73_72 202000.000000
Rwneg73_73 in73_73 sn73_73 202000.000000
Rwneg73_74 in73_74 sn73_74 202000.000000
Rwneg73_75 in73_75 sn73_75 202000.000000
Rwneg73_76 in73_76 sn73_76 202000.000000
Rwneg73_77 in73_77 sn73_77 202000.000000
Rwneg73_78 in73_78 sn73_78 202000.000000
Rwneg73_79 in73_79 sn73_79 78000.000000
Rwneg73_80 in73_80 sn73_80 78000.000000
Rwneg73_81 in73_81 sn73_81 78000.000000
Rwneg73_82 in73_82 sn73_82 78000.000000
Rwneg73_83 in73_83 sn73_83 202000.000000
Rwneg73_84 in73_84 sn73_84 202000.000000
Rwneg74_1 in74_1 sn74_1 202000.000000
Rwneg74_2 in74_2 sn74_2 202000.000000
Rwneg74_3 in74_3 sn74_3 202000.000000
Rwneg74_4 in74_4 sn74_4 78000.000000
Rwneg74_5 in74_5 sn74_5 78000.000000
Rwneg74_6 in74_6 sn74_6 202000.000000
Rwneg74_7 in74_7 sn74_7 202000.000000
Rwneg74_8 in74_8 sn74_8 78000.000000
Rwneg74_9 in74_9 sn74_9 78000.000000
Rwneg74_10 in74_10 sn74_10 202000.000000
Rwneg74_11 in74_11 sn74_11 78000.000000
Rwneg74_12 in74_12 sn74_12 78000.000000
Rwneg74_13 in74_13 sn74_13 78000.000000
Rwneg74_14 in74_14 sn74_14 202000.000000
Rwneg74_15 in74_15 sn74_15 78000.000000
Rwneg74_16 in74_16 sn74_16 78000.000000
Rwneg74_17 in74_17 sn74_17 78000.000000
Rwneg74_18 in74_18 sn74_18 78000.000000
Rwneg74_19 in74_19 sn74_19 78000.000000
Rwneg74_20 in74_20 sn74_20 202000.000000
Rwneg74_21 in74_21 sn74_21 202000.000000
Rwneg74_22 in74_22 sn74_22 78000.000000
Rwneg74_23 in74_23 sn74_23 202000.000000
Rwneg74_24 in74_24 sn74_24 202000.000000
Rwneg74_25 in74_25 sn74_25 202000.000000
Rwneg74_26 in74_26 sn74_26 78000.000000
Rwneg74_27 in74_27 sn74_27 78000.000000
Rwneg74_28 in74_28 sn74_28 78000.000000
Rwneg74_29 in74_29 sn74_29 78000.000000
Rwneg74_30 in74_30 sn74_30 202000.000000
Rwneg74_31 in74_31 sn74_31 78000.000000
Rwneg74_32 in74_32 sn74_32 202000.000000
Rwneg74_33 in74_33 sn74_33 78000.000000
Rwneg74_34 in74_34 sn74_34 202000.000000
Rwneg74_35 in74_35 sn74_35 78000.000000
Rwneg74_36 in74_36 sn74_36 202000.000000
Rwneg74_37 in74_37 sn74_37 202000.000000
Rwneg74_38 in74_38 sn74_38 202000.000000
Rwneg74_39 in74_39 sn74_39 78000.000000
Rwneg74_40 in74_40 sn74_40 202000.000000
Rwneg74_41 in74_41 sn74_41 202000.000000
Rwneg74_42 in74_42 sn74_42 202000.000000
Rwneg74_43 in74_43 sn74_43 202000.000000
Rwneg74_44 in74_44 sn74_44 78000.000000
Rwneg74_45 in74_45 sn74_45 78000.000000
Rwneg74_46 in74_46 sn74_46 202000.000000
Rwneg74_47 in74_47 sn74_47 202000.000000
Rwneg74_48 in74_48 sn74_48 202000.000000
Rwneg74_49 in74_49 sn74_49 202000.000000
Rwneg74_50 in74_50 sn74_50 202000.000000
Rwneg74_51 in74_51 sn74_51 202000.000000
Rwneg74_52 in74_52 sn74_52 202000.000000
Rwneg74_53 in74_53 sn74_53 202000.000000
Rwneg74_54 in74_54 sn74_54 78000.000000
Rwneg74_55 in74_55 sn74_55 78000.000000
Rwneg74_56 in74_56 sn74_56 202000.000000
Rwneg74_57 in74_57 sn74_57 78000.000000
Rwneg74_58 in74_58 sn74_58 78000.000000
Rwneg74_59 in74_59 sn74_59 202000.000000
Rwneg74_60 in74_60 sn74_60 202000.000000
Rwneg74_61 in74_61 sn74_61 78000.000000
Rwneg74_62 in74_62 sn74_62 202000.000000
Rwneg74_63 in74_63 sn74_63 202000.000000
Rwneg74_64 in74_64 sn74_64 78000.000000
Rwneg74_65 in74_65 sn74_65 78000.000000
Rwneg74_66 in74_66 sn74_66 202000.000000
Rwneg74_67 in74_67 sn74_67 78000.000000
Rwneg74_68 in74_68 sn74_68 78000.000000
Rwneg74_69 in74_69 sn74_69 202000.000000
Rwneg74_70 in74_70 sn74_70 78000.000000
Rwneg74_71 in74_71 sn74_71 202000.000000
Rwneg74_72 in74_72 sn74_72 78000.000000
Rwneg74_73 in74_73 sn74_73 202000.000000
Rwneg74_74 in74_74 sn74_74 78000.000000
Rwneg74_75 in74_75 sn74_75 78000.000000
Rwneg74_76 in74_76 sn74_76 202000.000000
Rwneg74_77 in74_77 sn74_77 78000.000000
Rwneg74_78 in74_78 sn74_78 202000.000000
Rwneg74_79 in74_79 sn74_79 202000.000000
Rwneg74_80 in74_80 sn74_80 78000.000000
Rwneg74_81 in74_81 sn74_81 202000.000000
Rwneg74_82 in74_82 sn74_82 202000.000000
Rwneg74_83 in74_83 sn74_83 202000.000000
Rwneg74_84 in74_84 sn74_84 202000.000000
Rwneg75_1 in75_1 sn75_1 202000.000000
Rwneg75_2 in75_2 sn75_2 78000.000000
Rwneg75_3 in75_3 sn75_3 78000.000000
Rwneg75_4 in75_4 sn75_4 78000.000000
Rwneg75_5 in75_5 sn75_5 78000.000000
Rwneg75_6 in75_6 sn75_6 78000.000000
Rwneg75_7 in75_7 sn75_7 202000.000000
Rwneg75_8 in75_8 sn75_8 202000.000000
Rwneg75_9 in75_9 sn75_9 202000.000000
Rwneg75_10 in75_10 sn75_10 202000.000000
Rwneg75_11 in75_11 sn75_11 78000.000000
Rwneg75_12 in75_12 sn75_12 202000.000000
Rwneg75_13 in75_13 sn75_13 78000.000000
Rwneg75_14 in75_14 sn75_14 202000.000000
Rwneg75_15 in75_15 sn75_15 78000.000000
Rwneg75_16 in75_16 sn75_16 78000.000000
Rwneg75_17 in75_17 sn75_17 202000.000000
Rwneg75_18 in75_18 sn75_18 78000.000000
Rwneg75_19 in75_19 sn75_19 78000.000000
Rwneg75_20 in75_20 sn75_20 78000.000000
Rwneg75_21 in75_21 sn75_21 78000.000000
Rwneg75_22 in75_22 sn75_22 202000.000000
Rwneg75_23 in75_23 sn75_23 202000.000000
Rwneg75_24 in75_24 sn75_24 78000.000000
Rwneg75_25 in75_25 sn75_25 78000.000000
Rwneg75_26 in75_26 sn75_26 202000.000000
Rwneg75_27 in75_27 sn75_27 202000.000000
Rwneg75_28 in75_28 sn75_28 78000.000000
Rwneg75_29 in75_29 sn75_29 78000.000000
Rwneg75_30 in75_30 sn75_30 78000.000000
Rwneg75_31 in75_31 sn75_31 202000.000000
Rwneg75_32 in75_32 sn75_32 202000.000000
Rwneg75_33 in75_33 sn75_33 78000.000000
Rwneg75_34 in75_34 sn75_34 202000.000000
Rwneg75_35 in75_35 sn75_35 202000.000000
Rwneg75_36 in75_36 sn75_36 78000.000000
Rwneg75_37 in75_37 sn75_37 202000.000000
Rwneg75_38 in75_38 sn75_38 78000.000000
Rwneg75_39 in75_39 sn75_39 78000.000000
Rwneg75_40 in75_40 sn75_40 78000.000000
Rwneg75_41 in75_41 sn75_41 202000.000000
Rwneg75_42 in75_42 sn75_42 202000.000000
Rwneg75_43 in75_43 sn75_43 78000.000000
Rwneg75_44 in75_44 sn75_44 78000.000000
Rwneg75_45 in75_45 sn75_45 78000.000000
Rwneg75_46 in75_46 sn75_46 202000.000000
Rwneg75_47 in75_47 sn75_47 78000.000000
Rwneg75_48 in75_48 sn75_48 78000.000000
Rwneg75_49 in75_49 sn75_49 202000.000000
Rwneg75_50 in75_50 sn75_50 78000.000000
Rwneg75_51 in75_51 sn75_51 202000.000000
Rwneg75_52 in75_52 sn75_52 78000.000000
Rwneg75_53 in75_53 sn75_53 78000.000000
Rwneg75_54 in75_54 sn75_54 78000.000000
Rwneg75_55 in75_55 sn75_55 78000.000000
Rwneg75_56 in75_56 sn75_56 202000.000000
Rwneg75_57 in75_57 sn75_57 78000.000000
Rwneg75_58 in75_58 sn75_58 202000.000000
Rwneg75_59 in75_59 sn75_59 202000.000000
Rwneg75_60 in75_60 sn75_60 202000.000000
Rwneg75_61 in75_61 sn75_61 202000.000000
Rwneg75_62 in75_62 sn75_62 202000.000000
Rwneg75_63 in75_63 sn75_63 202000.000000
Rwneg75_64 in75_64 sn75_64 202000.000000
Rwneg75_65 in75_65 sn75_65 78000.000000
Rwneg75_66 in75_66 sn75_66 202000.000000
Rwneg75_67 in75_67 sn75_67 78000.000000
Rwneg75_68 in75_68 sn75_68 202000.000000
Rwneg75_69 in75_69 sn75_69 202000.000000
Rwneg75_70 in75_70 sn75_70 78000.000000
Rwneg75_71 in75_71 sn75_71 78000.000000
Rwneg75_72 in75_72 sn75_72 202000.000000
Rwneg75_73 in75_73 sn75_73 202000.000000
Rwneg75_74 in75_74 sn75_74 202000.000000
Rwneg75_75 in75_75 sn75_75 78000.000000
Rwneg75_76 in75_76 sn75_76 202000.000000
Rwneg75_77 in75_77 sn75_77 78000.000000
Rwneg75_78 in75_78 sn75_78 202000.000000
Rwneg75_79 in75_79 sn75_79 202000.000000
Rwneg75_80 in75_80 sn75_80 202000.000000
Rwneg75_81 in75_81 sn75_81 78000.000000
Rwneg75_82 in75_82 sn75_82 202000.000000
Rwneg75_83 in75_83 sn75_83 78000.000000
Rwneg75_84 in75_84 sn75_84 78000.000000
Rwneg76_1 in76_1 sn76_1 78000.000000
Rwneg76_2 in76_2 sn76_2 202000.000000
Rwneg76_3 in76_3 sn76_3 78000.000000
Rwneg76_4 in76_4 sn76_4 78000.000000
Rwneg76_5 in76_5 sn76_5 202000.000000
Rwneg76_6 in76_6 sn76_6 78000.000000
Rwneg76_7 in76_7 sn76_7 202000.000000
Rwneg76_8 in76_8 sn76_8 78000.000000
Rwneg76_9 in76_9 sn76_9 78000.000000
Rwneg76_10 in76_10 sn76_10 202000.000000
Rwneg76_11 in76_11 sn76_11 202000.000000
Rwneg76_12 in76_12 sn76_12 78000.000000
Rwneg76_13 in76_13 sn76_13 78000.000000
Rwneg76_14 in76_14 sn76_14 78000.000000
Rwneg76_15 in76_15 sn76_15 202000.000000
Rwneg76_16 in76_16 sn76_16 78000.000000
Rwneg76_17 in76_17 sn76_17 202000.000000
Rwneg76_18 in76_18 sn76_18 78000.000000
Rwneg76_19 in76_19 sn76_19 202000.000000
Rwneg76_20 in76_20 sn76_20 202000.000000
Rwneg76_21 in76_21 sn76_21 78000.000000
Rwneg76_22 in76_22 sn76_22 78000.000000
Rwneg76_23 in76_23 sn76_23 78000.000000
Rwneg76_24 in76_24 sn76_24 202000.000000
Rwneg76_25 in76_25 sn76_25 202000.000000
Rwneg76_26 in76_26 sn76_26 78000.000000
Rwneg76_27 in76_27 sn76_27 78000.000000
Rwneg76_28 in76_28 sn76_28 202000.000000
Rwneg76_29 in76_29 sn76_29 78000.000000
Rwneg76_30 in76_30 sn76_30 202000.000000
Rwneg76_31 in76_31 sn76_31 78000.000000
Rwneg76_32 in76_32 sn76_32 202000.000000
Rwneg76_33 in76_33 sn76_33 202000.000000
Rwneg76_34 in76_34 sn76_34 202000.000000
Rwneg76_35 in76_35 sn76_35 78000.000000
Rwneg76_36 in76_36 sn76_36 202000.000000
Rwneg76_37 in76_37 sn76_37 202000.000000
Rwneg76_38 in76_38 sn76_38 78000.000000
Rwneg76_39 in76_39 sn76_39 78000.000000
Rwneg76_40 in76_40 sn76_40 78000.000000
Rwneg76_41 in76_41 sn76_41 78000.000000
Rwneg76_42 in76_42 sn76_42 202000.000000
Rwneg76_43 in76_43 sn76_43 78000.000000
Rwneg76_44 in76_44 sn76_44 202000.000000
Rwneg76_45 in76_45 sn76_45 78000.000000
Rwneg76_46 in76_46 sn76_46 202000.000000
Rwneg76_47 in76_47 sn76_47 202000.000000
Rwneg76_48 in76_48 sn76_48 78000.000000
Rwneg76_49 in76_49 sn76_49 202000.000000
Rwneg76_50 in76_50 sn76_50 202000.000000
Rwneg76_51 in76_51 sn76_51 202000.000000
Rwneg76_52 in76_52 sn76_52 202000.000000
Rwneg76_53 in76_53 sn76_53 202000.000000
Rwneg76_54 in76_54 sn76_54 202000.000000
Rwneg76_55 in76_55 sn76_55 202000.000000
Rwneg76_56 in76_56 sn76_56 202000.000000
Rwneg76_57 in76_57 sn76_57 78000.000000
Rwneg76_58 in76_58 sn76_58 78000.000000
Rwneg76_59 in76_59 sn76_59 78000.000000
Rwneg76_60 in76_60 sn76_60 202000.000000
Rwneg76_61 in76_61 sn76_61 202000.000000
Rwneg76_62 in76_62 sn76_62 202000.000000
Rwneg76_63 in76_63 sn76_63 78000.000000
Rwneg76_64 in76_64 sn76_64 202000.000000
Rwneg76_65 in76_65 sn76_65 78000.000000
Rwneg76_66 in76_66 sn76_66 202000.000000
Rwneg76_67 in76_67 sn76_67 78000.000000
Rwneg76_68 in76_68 sn76_68 78000.000000
Rwneg76_69 in76_69 sn76_69 202000.000000
Rwneg76_70 in76_70 sn76_70 78000.000000
Rwneg76_71 in76_71 sn76_71 78000.000000
Rwneg76_72 in76_72 sn76_72 78000.000000
Rwneg76_73 in76_73 sn76_73 78000.000000
Rwneg76_74 in76_74 sn76_74 78000.000000
Rwneg76_75 in76_75 sn76_75 78000.000000
Rwneg76_76 in76_76 sn76_76 202000.000000
Rwneg76_77 in76_77 sn76_77 78000.000000
Rwneg76_78 in76_78 sn76_78 202000.000000
Rwneg76_79 in76_79 sn76_79 202000.000000
Rwneg76_80 in76_80 sn76_80 202000.000000
Rwneg76_81 in76_81 sn76_81 202000.000000
Rwneg76_82 in76_82 sn76_82 202000.000000
Rwneg76_83 in76_83 sn76_83 78000.000000
Rwneg76_84 in76_84 sn76_84 78000.000000
Rwneg77_1 in77_1 sn77_1 202000.000000
Rwneg77_2 in77_2 sn77_2 202000.000000
Rwneg77_3 in77_3 sn77_3 202000.000000
Rwneg77_4 in77_4 sn77_4 202000.000000
Rwneg77_5 in77_5 sn77_5 202000.000000
Rwneg77_6 in77_6 sn77_6 78000.000000
Rwneg77_7 in77_7 sn77_7 202000.000000
Rwneg77_8 in77_8 sn77_8 202000.000000
Rwneg77_9 in77_9 sn77_9 78000.000000
Rwneg77_10 in77_10 sn77_10 202000.000000
Rwneg77_11 in77_11 sn77_11 202000.000000
Rwneg77_12 in77_12 sn77_12 202000.000000
Rwneg77_13 in77_13 sn77_13 202000.000000
Rwneg77_14 in77_14 sn77_14 202000.000000
Rwneg77_15 in77_15 sn77_15 202000.000000
Rwneg77_16 in77_16 sn77_16 78000.000000
Rwneg77_17 in77_17 sn77_17 202000.000000
Rwneg77_18 in77_18 sn77_18 78000.000000
Rwneg77_19 in77_19 sn77_19 78000.000000
Rwneg77_20 in77_20 sn77_20 78000.000000
Rwneg77_21 in77_21 sn77_21 78000.000000
Rwneg77_22 in77_22 sn77_22 78000.000000
Rwneg77_23 in77_23 sn77_23 78000.000000
Rwneg77_24 in77_24 sn77_24 78000.000000
Rwneg77_25 in77_25 sn77_25 202000.000000
Rwneg77_26 in77_26 sn77_26 78000.000000
Rwneg77_27 in77_27 sn77_27 202000.000000
Rwneg77_28 in77_28 sn77_28 202000.000000
Rwneg77_29 in77_29 sn77_29 202000.000000
Rwneg77_30 in77_30 sn77_30 202000.000000
Rwneg77_31 in77_31 sn77_31 202000.000000
Rwneg77_32 in77_32 sn77_32 202000.000000
Rwneg77_33 in77_33 sn77_33 78000.000000
Rwneg77_34 in77_34 sn77_34 202000.000000
Rwneg77_35 in77_35 sn77_35 202000.000000
Rwneg77_36 in77_36 sn77_36 202000.000000
Rwneg77_37 in77_37 sn77_37 78000.000000
Rwneg77_38 in77_38 sn77_38 78000.000000
Rwneg77_39 in77_39 sn77_39 202000.000000
Rwneg77_40 in77_40 sn77_40 78000.000000
Rwneg77_41 in77_41 sn77_41 78000.000000
Rwneg77_42 in77_42 sn77_42 202000.000000
Rwneg77_43 in77_43 sn77_43 78000.000000
Rwneg77_44 in77_44 sn77_44 202000.000000
Rwneg77_45 in77_45 sn77_45 78000.000000
Rwneg77_46 in77_46 sn77_46 202000.000000
Rwneg77_47 in77_47 sn77_47 202000.000000
Rwneg77_48 in77_48 sn77_48 78000.000000
Rwneg77_49 in77_49 sn77_49 202000.000000
Rwneg77_50 in77_50 sn77_50 202000.000000
Rwneg77_51 in77_51 sn77_51 78000.000000
Rwneg77_52 in77_52 sn77_52 78000.000000
Rwneg77_53 in77_53 sn77_53 78000.000000
Rwneg77_54 in77_54 sn77_54 78000.000000
Rwneg77_55 in77_55 sn77_55 78000.000000
Rwneg77_56 in77_56 sn77_56 78000.000000
Rwneg77_57 in77_57 sn77_57 78000.000000
Rwneg77_58 in77_58 sn77_58 202000.000000
Rwneg77_59 in77_59 sn77_59 202000.000000
Rwneg77_60 in77_60 sn77_60 78000.000000
Rwneg77_61 in77_61 sn77_61 78000.000000
Rwneg77_62 in77_62 sn77_62 202000.000000
Rwneg77_63 in77_63 sn77_63 78000.000000
Rwneg77_64 in77_64 sn77_64 78000.000000
Rwneg77_65 in77_65 sn77_65 78000.000000
Rwneg77_66 in77_66 sn77_66 78000.000000
Rwneg77_67 in77_67 sn77_67 202000.000000
Rwneg77_68 in77_68 sn77_68 202000.000000
Rwneg77_69 in77_69 sn77_69 202000.000000
Rwneg77_70 in77_70 sn77_70 78000.000000
Rwneg77_71 in77_71 sn77_71 78000.000000
Rwneg77_72 in77_72 sn77_72 78000.000000
Rwneg77_73 in77_73 sn77_73 78000.000000
Rwneg77_74 in77_74 sn77_74 202000.000000
Rwneg77_75 in77_75 sn77_75 202000.000000
Rwneg77_76 in77_76 sn77_76 202000.000000
Rwneg77_77 in77_77 sn77_77 78000.000000
Rwneg77_78 in77_78 sn77_78 78000.000000
Rwneg77_79 in77_79 sn77_79 78000.000000
Rwneg77_80 in77_80 sn77_80 202000.000000
Rwneg77_81 in77_81 sn77_81 202000.000000
Rwneg77_82 in77_82 sn77_82 78000.000000
Rwneg77_83 in77_83 sn77_83 78000.000000
Rwneg77_84 in77_84 sn77_84 78000.000000
Rwneg78_1 in78_1 sn78_1 202000.000000
Rwneg78_2 in78_2 sn78_2 202000.000000
Rwneg78_3 in78_3 sn78_3 202000.000000
Rwneg78_4 in78_4 sn78_4 202000.000000
Rwneg78_5 in78_5 sn78_5 202000.000000
Rwneg78_6 in78_6 sn78_6 202000.000000
Rwneg78_7 in78_7 sn78_7 202000.000000
Rwneg78_8 in78_8 sn78_8 78000.000000
Rwneg78_9 in78_9 sn78_9 78000.000000
Rwneg78_10 in78_10 sn78_10 202000.000000
Rwneg78_11 in78_11 sn78_11 78000.000000
Rwneg78_12 in78_12 sn78_12 78000.000000
Rwneg78_13 in78_13 sn78_13 202000.000000
Rwneg78_14 in78_14 sn78_14 202000.000000
Rwneg78_15 in78_15 sn78_15 202000.000000
Rwneg78_16 in78_16 sn78_16 78000.000000
Rwneg78_17 in78_17 sn78_17 202000.000000
Rwneg78_18 in78_18 sn78_18 78000.000000
Rwneg78_19 in78_19 sn78_19 202000.000000
Rwneg78_20 in78_20 sn78_20 202000.000000
Rwneg78_21 in78_21 sn78_21 78000.000000
Rwneg78_22 in78_22 sn78_22 78000.000000
Rwneg78_23 in78_23 sn78_23 78000.000000
Rwneg78_24 in78_24 sn78_24 202000.000000
Rwneg78_25 in78_25 sn78_25 78000.000000
Rwneg78_26 in78_26 sn78_26 202000.000000
Rwneg78_27 in78_27 sn78_27 78000.000000
Rwneg78_28 in78_28 sn78_28 78000.000000
Rwneg78_29 in78_29 sn78_29 78000.000000
Rwneg78_30 in78_30 sn78_30 202000.000000
Rwneg78_31 in78_31 sn78_31 78000.000000
Rwneg78_32 in78_32 sn78_32 78000.000000
Rwneg78_33 in78_33 sn78_33 202000.000000
Rwneg78_34 in78_34 sn78_34 78000.000000
Rwneg78_35 in78_35 sn78_35 78000.000000
Rwneg78_36 in78_36 sn78_36 78000.000000
Rwneg78_37 in78_37 sn78_37 78000.000000
Rwneg78_38 in78_38 sn78_38 202000.000000
Rwneg78_39 in78_39 sn78_39 202000.000000
Rwneg78_40 in78_40 sn78_40 78000.000000
Rwneg78_41 in78_41 sn78_41 78000.000000
Rwneg78_42 in78_42 sn78_42 202000.000000
Rwneg78_43 in78_43 sn78_43 78000.000000
Rwneg78_44 in78_44 sn78_44 202000.000000
Rwneg78_45 in78_45 sn78_45 78000.000000
Rwneg78_46 in78_46 sn78_46 202000.000000
Rwneg78_47 in78_47 sn78_47 202000.000000
Rwneg78_48 in78_48 sn78_48 202000.000000
Rwneg78_49 in78_49 sn78_49 202000.000000
Rwneg78_50 in78_50 sn78_50 202000.000000
Rwneg78_51 in78_51 sn78_51 202000.000000
Rwneg78_52 in78_52 sn78_52 202000.000000
Rwneg78_53 in78_53 sn78_53 78000.000000
Rwneg78_54 in78_54 sn78_54 202000.000000
Rwneg78_55 in78_55 sn78_55 78000.000000
Rwneg78_56 in78_56 sn78_56 78000.000000
Rwneg78_57 in78_57 sn78_57 202000.000000
Rwneg78_58 in78_58 sn78_58 78000.000000
Rwneg78_59 in78_59 sn78_59 202000.000000
Rwneg78_60 in78_60 sn78_60 202000.000000
Rwneg78_61 in78_61 sn78_61 78000.000000
Rwneg78_62 in78_62 sn78_62 202000.000000
Rwneg78_63 in78_63 sn78_63 202000.000000
Rwneg78_64 in78_64 sn78_64 202000.000000
Rwneg78_65 in78_65 sn78_65 78000.000000
Rwneg78_66 in78_66 sn78_66 78000.000000
Rwneg78_67 in78_67 sn78_67 202000.000000
Rwneg78_68 in78_68 sn78_68 78000.000000
Rwneg78_69 in78_69 sn78_69 78000.000000
Rwneg78_70 in78_70 sn78_70 78000.000000
Rwneg78_71 in78_71 sn78_71 78000.000000
Rwneg78_72 in78_72 sn78_72 202000.000000
Rwneg78_73 in78_73 sn78_73 78000.000000
Rwneg78_74 in78_74 sn78_74 202000.000000
Rwneg78_75 in78_75 sn78_75 202000.000000
Rwneg78_76 in78_76 sn78_76 78000.000000
Rwneg78_77 in78_77 sn78_77 78000.000000
Rwneg78_78 in78_78 sn78_78 78000.000000
Rwneg78_79 in78_79 sn78_79 78000.000000
Rwneg78_80 in78_80 sn78_80 78000.000000
Rwneg78_81 in78_81 sn78_81 202000.000000
Rwneg78_82 in78_82 sn78_82 78000.000000
Rwneg78_83 in78_83 sn78_83 202000.000000
Rwneg78_84 in78_84 sn78_84 202000.000000
Rwneg79_1 in79_1 sn79_1 78000.000000
Rwneg79_2 in79_2 sn79_2 78000.000000
Rwneg79_3 in79_3 sn79_3 202000.000000
Rwneg79_4 in79_4 sn79_4 202000.000000
Rwneg79_5 in79_5 sn79_5 202000.000000
Rwneg79_6 in79_6 sn79_6 78000.000000
Rwneg79_7 in79_7 sn79_7 78000.000000
Rwneg79_8 in79_8 sn79_8 202000.000000
Rwneg79_9 in79_9 sn79_9 202000.000000
Rwneg79_10 in79_10 sn79_10 78000.000000
Rwneg79_11 in79_11 sn79_11 202000.000000
Rwneg79_12 in79_12 sn79_12 78000.000000
Rwneg79_13 in79_13 sn79_13 78000.000000
Rwneg79_14 in79_14 sn79_14 78000.000000
Rwneg79_15 in79_15 sn79_15 202000.000000
Rwneg79_16 in79_16 sn79_16 78000.000000
Rwneg79_17 in79_17 sn79_17 78000.000000
Rwneg79_18 in79_18 sn79_18 202000.000000
Rwneg79_19 in79_19 sn79_19 78000.000000
Rwneg79_20 in79_20 sn79_20 202000.000000
Rwneg79_21 in79_21 sn79_21 78000.000000
Rwneg79_22 in79_22 sn79_22 202000.000000
Rwneg79_23 in79_23 sn79_23 78000.000000
Rwneg79_24 in79_24 sn79_24 78000.000000
Rwneg79_25 in79_25 sn79_25 202000.000000
Rwneg79_26 in79_26 sn79_26 202000.000000
Rwneg79_27 in79_27 sn79_27 78000.000000
Rwneg79_28 in79_28 sn79_28 202000.000000
Rwneg79_29 in79_29 sn79_29 78000.000000
Rwneg79_30 in79_30 sn79_30 78000.000000
Rwneg79_31 in79_31 sn79_31 78000.000000
Rwneg79_32 in79_32 sn79_32 78000.000000
Rwneg79_33 in79_33 sn79_33 202000.000000
Rwneg79_34 in79_34 sn79_34 78000.000000
Rwneg79_35 in79_35 sn79_35 202000.000000
Rwneg79_36 in79_36 sn79_36 78000.000000
Rwneg79_37 in79_37 sn79_37 202000.000000
Rwneg79_38 in79_38 sn79_38 78000.000000
Rwneg79_39 in79_39 sn79_39 78000.000000
Rwneg79_40 in79_40 sn79_40 78000.000000
Rwneg79_41 in79_41 sn79_41 78000.000000
Rwneg79_42 in79_42 sn79_42 202000.000000
Rwneg79_43 in79_43 sn79_43 202000.000000
Rwneg79_44 in79_44 sn79_44 78000.000000
Rwneg79_45 in79_45 sn79_45 202000.000000
Rwneg79_46 in79_46 sn79_46 202000.000000
Rwneg79_47 in79_47 sn79_47 78000.000000
Rwneg79_48 in79_48 sn79_48 78000.000000
Rwneg79_49 in79_49 sn79_49 202000.000000
Rwneg79_50 in79_50 sn79_50 202000.000000
Rwneg79_51 in79_51 sn79_51 202000.000000
Rwneg79_52 in79_52 sn79_52 202000.000000
Rwneg79_53 in79_53 sn79_53 78000.000000
Rwneg79_54 in79_54 sn79_54 202000.000000
Rwneg79_55 in79_55 sn79_55 202000.000000
Rwneg79_56 in79_56 sn79_56 78000.000000
Rwneg79_57 in79_57 sn79_57 202000.000000
Rwneg79_58 in79_58 sn79_58 78000.000000
Rwneg79_59 in79_59 sn79_59 202000.000000
Rwneg79_60 in79_60 sn79_60 78000.000000
Rwneg79_61 in79_61 sn79_61 202000.000000
Rwneg79_62 in79_62 sn79_62 78000.000000
Rwneg79_63 in79_63 sn79_63 78000.000000
Rwneg79_64 in79_64 sn79_64 78000.000000
Rwneg79_65 in79_65 sn79_65 78000.000000
Rwneg79_66 in79_66 sn79_66 78000.000000
Rwneg79_67 in79_67 sn79_67 78000.000000
Rwneg79_68 in79_68 sn79_68 78000.000000
Rwneg79_69 in79_69 sn79_69 202000.000000
Rwneg79_70 in79_70 sn79_70 78000.000000
Rwneg79_71 in79_71 sn79_71 202000.000000
Rwneg79_72 in79_72 sn79_72 202000.000000
Rwneg79_73 in79_73 sn79_73 202000.000000
Rwneg79_74 in79_74 sn79_74 202000.000000
Rwneg79_75 in79_75 sn79_75 202000.000000
Rwneg79_76 in79_76 sn79_76 78000.000000
Rwneg79_77 in79_77 sn79_77 78000.000000
Rwneg79_78 in79_78 sn79_78 202000.000000
Rwneg79_79 in79_79 sn79_79 78000.000000
Rwneg79_80 in79_80 sn79_80 202000.000000
Rwneg79_81 in79_81 sn79_81 78000.000000
Rwneg79_82 in79_82 sn79_82 78000.000000
Rwneg79_83 in79_83 sn79_83 78000.000000
Rwneg79_84 in79_84 sn79_84 202000.000000
Rwneg80_1 in80_1 sn80_1 202000.000000
Rwneg80_2 in80_2 sn80_2 78000.000000
Rwneg80_3 in80_3 sn80_3 202000.000000
Rwneg80_4 in80_4 sn80_4 202000.000000
Rwneg80_5 in80_5 sn80_5 202000.000000
Rwneg80_6 in80_6 sn80_6 78000.000000
Rwneg80_7 in80_7 sn80_7 78000.000000
Rwneg80_8 in80_8 sn80_8 202000.000000
Rwneg80_9 in80_9 sn80_9 202000.000000
Rwneg80_10 in80_10 sn80_10 202000.000000
Rwneg80_11 in80_11 sn80_11 78000.000000
Rwneg80_12 in80_12 sn80_12 202000.000000
Rwneg80_13 in80_13 sn80_13 202000.000000
Rwneg80_14 in80_14 sn80_14 202000.000000
Rwneg80_15 in80_15 sn80_15 78000.000000
Rwneg80_16 in80_16 sn80_16 78000.000000
Rwneg80_17 in80_17 sn80_17 78000.000000
Rwneg80_18 in80_18 sn80_18 78000.000000
Rwneg80_19 in80_19 sn80_19 202000.000000
Rwneg80_20 in80_20 sn80_20 202000.000000
Rwneg80_21 in80_21 sn80_21 202000.000000
Rwneg80_22 in80_22 sn80_22 202000.000000
Rwneg80_23 in80_23 sn80_23 202000.000000
Rwneg80_24 in80_24 sn80_24 78000.000000
Rwneg80_25 in80_25 sn80_25 202000.000000
Rwneg80_26 in80_26 sn80_26 202000.000000
Rwneg80_27 in80_27 sn80_27 202000.000000
Rwneg80_28 in80_28 sn80_28 202000.000000
Rwneg80_29 in80_29 sn80_29 78000.000000
Rwneg80_30 in80_30 sn80_30 202000.000000
Rwneg80_31 in80_31 sn80_31 78000.000000
Rwneg80_32 in80_32 sn80_32 202000.000000
Rwneg80_33 in80_33 sn80_33 78000.000000
Rwneg80_34 in80_34 sn80_34 202000.000000
Rwneg80_35 in80_35 sn80_35 202000.000000
Rwneg80_36 in80_36 sn80_36 202000.000000
Rwneg80_37 in80_37 sn80_37 202000.000000
Rwneg80_38 in80_38 sn80_38 202000.000000
Rwneg80_39 in80_39 sn80_39 202000.000000
Rwneg80_40 in80_40 sn80_40 202000.000000
Rwneg80_41 in80_41 sn80_41 78000.000000
Rwneg80_42 in80_42 sn80_42 78000.000000
Rwneg80_43 in80_43 sn80_43 202000.000000
Rwneg80_44 in80_44 sn80_44 202000.000000
Rwneg80_45 in80_45 sn80_45 202000.000000
Rwneg80_46 in80_46 sn80_46 78000.000000
Rwneg80_47 in80_47 sn80_47 78000.000000
Rwneg80_48 in80_48 sn80_48 202000.000000
Rwneg80_49 in80_49 sn80_49 202000.000000
Rwneg80_50 in80_50 sn80_50 202000.000000
Rwneg80_51 in80_51 sn80_51 202000.000000
Rwneg80_52 in80_52 sn80_52 202000.000000
Rwneg80_53 in80_53 sn80_53 78000.000000
Rwneg80_54 in80_54 sn80_54 202000.000000
Rwneg80_55 in80_55 sn80_55 202000.000000
Rwneg80_56 in80_56 sn80_56 202000.000000
Rwneg80_57 in80_57 sn80_57 202000.000000
Rwneg80_58 in80_58 sn80_58 78000.000000
Rwneg80_59 in80_59 sn80_59 202000.000000
Rwneg80_60 in80_60 sn80_60 202000.000000
Rwneg80_61 in80_61 sn80_61 202000.000000
Rwneg80_62 in80_62 sn80_62 78000.000000
Rwneg80_63 in80_63 sn80_63 202000.000000
Rwneg80_64 in80_64 sn80_64 78000.000000
Rwneg80_65 in80_65 sn80_65 78000.000000
Rwneg80_66 in80_66 sn80_66 202000.000000
Rwneg80_67 in80_67 sn80_67 202000.000000
Rwneg80_68 in80_68 sn80_68 78000.000000
Rwneg80_69 in80_69 sn80_69 78000.000000
Rwneg80_70 in80_70 sn80_70 202000.000000
Rwneg80_71 in80_71 sn80_71 202000.000000
Rwneg80_72 in80_72 sn80_72 202000.000000
Rwneg80_73 in80_73 sn80_73 202000.000000
Rwneg80_74 in80_74 sn80_74 202000.000000
Rwneg80_75 in80_75 sn80_75 202000.000000
Rwneg80_76 in80_76 sn80_76 202000.000000
Rwneg80_77 in80_77 sn80_77 78000.000000
Rwneg80_78 in80_78 sn80_78 78000.000000
Rwneg80_79 in80_79 sn80_79 202000.000000
Rwneg80_80 in80_80 sn80_80 202000.000000
Rwneg80_81 in80_81 sn80_81 78000.000000
Rwneg80_82 in80_82 sn80_82 202000.000000
Rwneg80_83 in80_83 sn80_83 78000.000000
Rwneg80_84 in80_84 sn80_84 78000.000000
Rwneg81_1 in81_1 sn81_1 202000.000000
Rwneg81_2 in81_2 sn81_2 202000.000000
Rwneg81_3 in81_3 sn81_3 202000.000000
Rwneg81_4 in81_4 sn81_4 202000.000000
Rwneg81_5 in81_5 sn81_5 202000.000000
Rwneg81_6 in81_6 sn81_6 78000.000000
Rwneg81_7 in81_7 sn81_7 202000.000000
Rwneg81_8 in81_8 sn81_8 202000.000000
Rwneg81_9 in81_9 sn81_9 78000.000000
Rwneg81_10 in81_10 sn81_10 202000.000000
Rwneg81_11 in81_11 sn81_11 202000.000000
Rwneg81_12 in81_12 sn81_12 78000.000000
Rwneg81_13 in81_13 sn81_13 78000.000000
Rwneg81_14 in81_14 sn81_14 202000.000000
Rwneg81_15 in81_15 sn81_15 202000.000000
Rwneg81_16 in81_16 sn81_16 202000.000000
Rwneg81_17 in81_17 sn81_17 78000.000000
Rwneg81_18 in81_18 sn81_18 202000.000000
Rwneg81_19 in81_19 sn81_19 202000.000000
Rwneg81_20 in81_20 sn81_20 202000.000000
Rwneg81_21 in81_21 sn81_21 78000.000000
Rwneg81_22 in81_22 sn81_22 78000.000000
Rwneg81_23 in81_23 sn81_23 202000.000000
Rwneg81_24 in81_24 sn81_24 78000.000000
Rwneg81_25 in81_25 sn81_25 78000.000000
Rwneg81_26 in81_26 sn81_26 78000.000000
Rwneg81_27 in81_27 sn81_27 202000.000000
Rwneg81_28 in81_28 sn81_28 202000.000000
Rwneg81_29 in81_29 sn81_29 78000.000000
Rwneg81_30 in81_30 sn81_30 78000.000000
Rwneg81_31 in81_31 sn81_31 202000.000000
Rwneg81_32 in81_32 sn81_32 202000.000000
Rwneg81_33 in81_33 sn81_33 202000.000000
Rwneg81_34 in81_34 sn81_34 78000.000000
Rwneg81_35 in81_35 sn81_35 202000.000000
Rwneg81_36 in81_36 sn81_36 78000.000000
Rwneg81_37 in81_37 sn81_37 78000.000000
Rwneg81_38 in81_38 sn81_38 78000.000000
Rwneg81_39 in81_39 sn81_39 202000.000000
Rwneg81_40 in81_40 sn81_40 78000.000000
Rwneg81_41 in81_41 sn81_41 78000.000000
Rwneg81_42 in81_42 sn81_42 202000.000000
Rwneg81_43 in81_43 sn81_43 202000.000000
Rwneg81_44 in81_44 sn81_44 78000.000000
Rwneg81_45 in81_45 sn81_45 202000.000000
Rwneg81_46 in81_46 sn81_46 78000.000000
Rwneg81_47 in81_47 sn81_47 78000.000000
Rwneg81_48 in81_48 sn81_48 78000.000000
Rwneg81_49 in81_49 sn81_49 202000.000000
Rwneg81_50 in81_50 sn81_50 202000.000000
Rwneg81_51 in81_51 sn81_51 202000.000000
Rwneg81_52 in81_52 sn81_52 202000.000000
Rwneg81_53 in81_53 sn81_53 202000.000000
Rwneg81_54 in81_54 sn81_54 202000.000000
Rwneg81_55 in81_55 sn81_55 78000.000000
Rwneg81_56 in81_56 sn81_56 78000.000000
Rwneg81_57 in81_57 sn81_57 78000.000000
Rwneg81_58 in81_58 sn81_58 202000.000000
Rwneg81_59 in81_59 sn81_59 78000.000000
Rwneg81_60 in81_60 sn81_60 202000.000000
Rwneg81_61 in81_61 sn81_61 78000.000000
Rwneg81_62 in81_62 sn81_62 78000.000000
Rwneg81_63 in81_63 sn81_63 78000.000000
Rwneg81_64 in81_64 sn81_64 202000.000000
Rwneg81_65 in81_65 sn81_65 78000.000000
Rwneg81_66 in81_66 sn81_66 202000.000000
Rwneg81_67 in81_67 sn81_67 78000.000000
Rwneg81_68 in81_68 sn81_68 78000.000000
Rwneg81_69 in81_69 sn81_69 202000.000000
Rwneg81_70 in81_70 sn81_70 202000.000000
Rwneg81_71 in81_71 sn81_71 78000.000000
Rwneg81_72 in81_72 sn81_72 202000.000000
Rwneg81_73 in81_73 sn81_73 78000.000000
Rwneg81_74 in81_74 sn81_74 78000.000000
Rwneg81_75 in81_75 sn81_75 202000.000000
Rwneg81_76 in81_76 sn81_76 78000.000000
Rwneg81_77 in81_77 sn81_77 78000.000000
Rwneg81_78 in81_78 sn81_78 78000.000000
Rwneg81_79 in81_79 sn81_79 78000.000000
Rwneg81_80 in81_80 sn81_80 202000.000000
Rwneg81_81 in81_81 sn81_81 202000.000000
Rwneg81_82 in81_82 sn81_82 78000.000000
Rwneg81_83 in81_83 sn81_83 202000.000000
Rwneg81_84 in81_84 sn81_84 202000.000000
Rwneg82_1 in82_1 sn82_1 78000.000000
Rwneg82_2 in82_2 sn82_2 78000.000000
Rwneg82_3 in82_3 sn82_3 78000.000000
Rwneg82_4 in82_4 sn82_4 202000.000000
Rwneg82_5 in82_5 sn82_5 202000.000000
Rwneg82_6 in82_6 sn82_6 78000.000000
Rwneg82_7 in82_7 sn82_7 78000.000000
Rwneg82_8 in82_8 sn82_8 202000.000000
Rwneg82_9 in82_9 sn82_9 202000.000000
Rwneg82_10 in82_10 sn82_10 78000.000000
Rwneg82_11 in82_11 sn82_11 202000.000000
Rwneg82_12 in82_12 sn82_12 202000.000000
Rwneg82_13 in82_13 sn82_13 202000.000000
Rwneg82_14 in82_14 sn82_14 78000.000000
Rwneg82_15 in82_15 sn82_15 202000.000000
Rwneg82_16 in82_16 sn82_16 202000.000000
Rwneg82_17 in82_17 sn82_17 78000.000000
Rwneg82_18 in82_18 sn82_18 202000.000000
Rwneg82_19 in82_19 sn82_19 202000.000000
Rwneg82_20 in82_20 sn82_20 202000.000000
Rwneg82_21 in82_21 sn82_21 202000.000000
Rwneg82_22 in82_22 sn82_22 202000.000000
Rwneg82_23 in82_23 sn82_23 202000.000000
Rwneg82_24 in82_24 sn82_24 202000.000000
Rwneg82_25 in82_25 sn82_25 78000.000000
Rwneg82_26 in82_26 sn82_26 78000.000000
Rwneg82_27 in82_27 sn82_27 202000.000000
Rwneg82_28 in82_28 sn82_28 202000.000000
Rwneg82_29 in82_29 sn82_29 78000.000000
Rwneg82_30 in82_30 sn82_30 202000.000000
Rwneg82_31 in82_31 sn82_31 78000.000000
Rwneg82_32 in82_32 sn82_32 78000.000000
Rwneg82_33 in82_33 sn82_33 202000.000000
Rwneg82_34 in82_34 sn82_34 78000.000000
Rwneg82_35 in82_35 sn82_35 202000.000000
Rwneg82_36 in82_36 sn82_36 78000.000000
Rwneg82_37 in82_37 sn82_37 78000.000000
Rwneg82_38 in82_38 sn82_38 78000.000000
Rwneg82_39 in82_39 sn82_39 202000.000000
Rwneg82_40 in82_40 sn82_40 78000.000000
Rwneg82_41 in82_41 sn82_41 202000.000000
Rwneg82_42 in82_42 sn82_42 78000.000000
Rwneg82_43 in82_43 sn82_43 202000.000000
Rwneg82_44 in82_44 sn82_44 78000.000000
Rwneg82_45 in82_45 sn82_45 202000.000000
Rwneg82_46 in82_46 sn82_46 78000.000000
Rwneg82_47 in82_47 sn82_47 78000.000000
Rwneg82_48 in82_48 sn82_48 202000.000000
Rwneg82_49 in82_49 sn82_49 202000.000000
Rwneg82_50 in82_50 sn82_50 78000.000000
Rwneg82_51 in82_51 sn82_51 202000.000000
Rwneg82_52 in82_52 sn82_52 78000.000000
Rwneg82_53 in82_53 sn82_53 78000.000000
Rwneg82_54 in82_54 sn82_54 78000.000000
Rwneg82_55 in82_55 sn82_55 202000.000000
Rwneg82_56 in82_56 sn82_56 202000.000000
Rwneg82_57 in82_57 sn82_57 202000.000000
Rwneg82_58 in82_58 sn82_58 78000.000000
Rwneg82_59 in82_59 sn82_59 78000.000000
Rwneg82_60 in82_60 sn82_60 78000.000000
Rwneg82_61 in82_61 sn82_61 202000.000000
Rwneg82_62 in82_62 sn82_62 202000.000000
Rwneg82_63 in82_63 sn82_63 202000.000000
Rwneg82_64 in82_64 sn82_64 78000.000000
Rwneg82_65 in82_65 sn82_65 202000.000000
Rwneg82_66 in82_66 sn82_66 202000.000000
Rwneg82_67 in82_67 sn82_67 78000.000000
Rwneg82_68 in82_68 sn82_68 202000.000000
Rwneg82_69 in82_69 sn82_69 202000.000000
Rwneg82_70 in82_70 sn82_70 202000.000000
Rwneg82_71 in82_71 sn82_71 202000.000000
Rwneg82_72 in82_72 sn82_72 78000.000000
Rwneg82_73 in82_73 sn82_73 202000.000000
Rwneg82_74 in82_74 sn82_74 78000.000000
Rwneg82_75 in82_75 sn82_75 78000.000000
Rwneg82_76 in82_76 sn82_76 78000.000000
Rwneg82_77 in82_77 sn82_77 78000.000000
Rwneg82_78 in82_78 sn82_78 78000.000000
Rwneg82_79 in82_79 sn82_79 78000.000000
Rwneg82_80 in82_80 sn82_80 202000.000000
Rwneg82_81 in82_81 sn82_81 202000.000000
Rwneg82_82 in82_82 sn82_82 202000.000000
Rwneg82_83 in82_83 sn82_83 202000.000000
Rwneg82_84 in82_84 sn82_84 202000.000000
Rwneg83_1 in83_1 sn83_1 202000.000000
Rwneg83_2 in83_2 sn83_2 202000.000000
Rwneg83_3 in83_3 sn83_3 78000.000000
Rwneg83_4 in83_4 sn83_4 202000.000000
Rwneg83_5 in83_5 sn83_5 202000.000000
Rwneg83_6 in83_6 sn83_6 78000.000000
Rwneg83_7 in83_7 sn83_7 202000.000000
Rwneg83_8 in83_8 sn83_8 202000.000000
Rwneg83_9 in83_9 sn83_9 202000.000000
Rwneg83_10 in83_10 sn83_10 78000.000000
Rwneg83_11 in83_11 sn83_11 78000.000000
Rwneg83_12 in83_12 sn83_12 202000.000000
Rwneg83_13 in83_13 sn83_13 78000.000000
Rwneg83_14 in83_14 sn83_14 78000.000000
Rwneg83_15 in83_15 sn83_15 78000.000000
Rwneg83_16 in83_16 sn83_16 202000.000000
Rwneg83_17 in83_17 sn83_17 202000.000000
Rwneg83_18 in83_18 sn83_18 202000.000000
Rwneg83_19 in83_19 sn83_19 202000.000000
Rwneg83_20 in83_20 sn83_20 202000.000000
Rwneg83_21 in83_21 sn83_21 202000.000000
Rwneg83_22 in83_22 sn83_22 202000.000000
Rwneg83_23 in83_23 sn83_23 78000.000000
Rwneg83_24 in83_24 sn83_24 202000.000000
Rwneg83_25 in83_25 sn83_25 202000.000000
Rwneg83_26 in83_26 sn83_26 202000.000000
Rwneg83_27 in83_27 sn83_27 202000.000000
Rwneg83_28 in83_28 sn83_28 78000.000000
Rwneg83_29 in83_29 sn83_29 78000.000000
Rwneg83_30 in83_30 sn83_30 78000.000000
Rwneg83_31 in83_31 sn83_31 78000.000000
Rwneg83_32 in83_32 sn83_32 202000.000000
Rwneg83_33 in83_33 sn83_33 202000.000000
Rwneg83_34 in83_34 sn83_34 78000.000000
Rwneg83_35 in83_35 sn83_35 78000.000000
Rwneg83_36 in83_36 sn83_36 78000.000000
Rwneg83_37 in83_37 sn83_37 202000.000000
Rwneg83_38 in83_38 sn83_38 78000.000000
Rwneg83_39 in83_39 sn83_39 78000.000000
Rwneg83_40 in83_40 sn83_40 78000.000000
Rwneg83_41 in83_41 sn83_41 78000.000000
Rwneg83_42 in83_42 sn83_42 202000.000000
Rwneg83_43 in83_43 sn83_43 202000.000000
Rwneg83_44 in83_44 sn83_44 202000.000000
Rwneg83_45 in83_45 sn83_45 78000.000000
Rwneg83_46 in83_46 sn83_46 78000.000000
Rwneg83_47 in83_47 sn83_47 78000.000000
Rwneg83_48 in83_48 sn83_48 202000.000000
Rwneg83_49 in83_49 sn83_49 78000.000000
Rwneg83_50 in83_50 sn83_50 78000.000000
Rwneg83_51 in83_51 sn83_51 78000.000000
Rwneg83_52 in83_52 sn83_52 202000.000000
Rwneg83_53 in83_53 sn83_53 78000.000000
Rwneg83_54 in83_54 sn83_54 202000.000000
Rwneg83_55 in83_55 sn83_55 78000.000000
Rwneg83_56 in83_56 sn83_56 78000.000000
Rwneg83_57 in83_57 sn83_57 78000.000000
Rwneg83_58 in83_58 sn83_58 78000.000000
Rwneg83_59 in83_59 sn83_59 202000.000000
Rwneg83_60 in83_60 sn83_60 202000.000000
Rwneg83_61 in83_61 sn83_61 78000.000000
Rwneg83_62 in83_62 sn83_62 202000.000000
Rwneg83_63 in83_63 sn83_63 202000.000000
Rwneg83_64 in83_64 sn83_64 202000.000000
Rwneg83_65 in83_65 sn83_65 202000.000000
Rwneg83_66 in83_66 sn83_66 202000.000000
Rwneg83_67 in83_67 sn83_67 78000.000000
Rwneg83_68 in83_68 sn83_68 78000.000000
Rwneg83_69 in83_69 sn83_69 202000.000000
Rwneg83_70 in83_70 sn83_70 78000.000000
Rwneg83_71 in83_71 sn83_71 78000.000000
Rwneg83_72 in83_72 sn83_72 78000.000000
Rwneg83_73 in83_73 sn83_73 78000.000000
Rwneg83_74 in83_74 sn83_74 78000.000000
Rwneg83_75 in83_75 sn83_75 78000.000000
Rwneg83_76 in83_76 sn83_76 78000.000000
Rwneg83_77 in83_77 sn83_77 78000.000000
Rwneg83_78 in83_78 sn83_78 78000.000000
Rwneg83_79 in83_79 sn83_79 78000.000000
Rwneg83_80 in83_80 sn83_80 202000.000000
Rwneg83_81 in83_81 sn83_81 202000.000000
Rwneg83_82 in83_82 sn83_82 202000.000000
Rwneg83_83 in83_83 sn83_83 202000.000000
Rwneg83_84 in83_84 sn83_84 202000.000000
Rwneg84_1 in84_1 sn84_1 78000.000000
Rwneg84_2 in84_2 sn84_2 78000.000000
Rwneg84_3 in84_3 sn84_3 78000.000000
Rwneg84_4 in84_4 sn84_4 78000.000000
Rwneg84_5 in84_5 sn84_5 78000.000000
Rwneg84_6 in84_6 sn84_6 78000.000000
Rwneg84_7 in84_7 sn84_7 78000.000000
Rwneg84_8 in84_8 sn84_8 202000.000000
Rwneg84_9 in84_9 sn84_9 202000.000000
Rwneg84_10 in84_10 sn84_10 78000.000000
Rwneg84_11 in84_11 sn84_11 202000.000000
Rwneg84_12 in84_12 sn84_12 202000.000000
Rwneg84_13 in84_13 sn84_13 78000.000000
Rwneg84_14 in84_14 sn84_14 78000.000000
Rwneg84_15 in84_15 sn84_15 78000.000000
Rwneg84_16 in84_16 sn84_16 202000.000000
Rwneg84_17 in84_17 sn84_17 202000.000000
Rwneg84_18 in84_18 sn84_18 202000.000000
Rwneg84_19 in84_19 sn84_19 78000.000000
Rwneg84_20 in84_20 sn84_20 78000.000000
Rwneg84_21 in84_21 sn84_21 202000.000000
Rwneg84_22 in84_22 sn84_22 202000.000000
Rwneg84_23 in84_23 sn84_23 202000.000000
Rwneg84_24 in84_24 sn84_24 202000.000000
Rwneg84_25 in84_25 sn84_25 78000.000000
Rwneg84_26 in84_26 sn84_26 202000.000000
Rwneg84_27 in84_27 sn84_27 202000.000000
Rwneg84_28 in84_28 sn84_28 202000.000000
Rwneg84_29 in84_29 sn84_29 78000.000000
Rwneg84_30 in84_30 sn84_30 202000.000000
Rwneg84_31 in84_31 sn84_31 202000.000000
Rwneg84_32 in84_32 sn84_32 202000.000000
Rwneg84_33 in84_33 sn84_33 78000.000000
Rwneg84_34 in84_34 sn84_34 202000.000000
Rwneg84_35 in84_35 sn84_35 78000.000000
Rwneg84_36 in84_36 sn84_36 202000.000000
Rwneg84_37 in84_37 sn84_37 202000.000000
Rwneg84_38 in84_38 sn84_38 78000.000000
Rwneg84_39 in84_39 sn84_39 78000.000000
Rwneg84_40 in84_40 sn84_40 202000.000000
Rwneg84_41 in84_41 sn84_41 202000.000000
Rwneg84_42 in84_42 sn84_42 78000.000000
Rwneg84_43 in84_43 sn84_43 202000.000000
Rwneg84_44 in84_44 sn84_44 78000.000000
Rwneg84_45 in84_45 sn84_45 78000.000000
Rwneg84_46 in84_46 sn84_46 78000.000000
Rwneg84_47 in84_47 sn84_47 78000.000000
Rwneg84_48 in84_48 sn84_48 202000.000000
Rwneg84_49 in84_49 sn84_49 78000.000000
Rwneg84_50 in84_50 sn84_50 78000.000000
Rwneg84_51 in84_51 sn84_51 202000.000000
Rwneg84_52 in84_52 sn84_52 202000.000000
Rwneg84_53 in84_53 sn84_53 202000.000000
Rwneg84_54 in84_54 sn84_54 202000.000000
Rwneg84_55 in84_55 sn84_55 78000.000000
Rwneg84_56 in84_56 sn84_56 202000.000000
Rwneg84_57 in84_57 sn84_57 202000.000000
Rwneg84_58 in84_58 sn84_58 202000.000000
Rwneg84_59 in84_59 sn84_59 78000.000000
Rwneg84_60 in84_60 sn84_60 78000.000000
Rwneg84_61 in84_61 sn84_61 202000.000000
Rwneg84_62 in84_62 sn84_62 78000.000000
Rwneg84_63 in84_63 sn84_63 78000.000000
Rwneg84_64 in84_64 sn84_64 202000.000000
Rwneg84_65 in84_65 sn84_65 202000.000000
Rwneg84_66 in84_66 sn84_66 202000.000000
Rwneg84_67 in84_67 sn84_67 202000.000000
Rwneg84_68 in84_68 sn84_68 202000.000000
Rwneg84_69 in84_69 sn84_69 202000.000000
Rwneg84_70 in84_70 sn84_70 78000.000000
Rwneg84_71 in84_71 sn84_71 202000.000000
Rwneg84_72 in84_72 sn84_72 78000.000000
Rwneg84_73 in84_73 sn84_73 202000.000000
Rwneg84_74 in84_74 sn84_74 202000.000000
Rwneg84_75 in84_75 sn84_75 78000.000000
Rwneg84_76 in84_76 sn84_76 202000.000000
Rwneg84_77 in84_77 sn84_77 78000.000000
Rwneg84_78 in84_78 sn84_78 202000.000000
Rwneg84_79 in84_79 sn84_79 202000.000000
Rwneg84_80 in84_80 sn84_80 202000.000000
Rwneg84_81 in84_81 sn84_81 78000.000000
Rwneg84_82 in84_82 sn84_82 202000.000000
Rwneg84_83 in84_83 sn84_83 78000.000000
Rwneg84_84 in84_84 sn84_84 78000.000000
Rwneg85_1 in85_1 sn85_1 78000.000000
Rwneg85_2 in85_2 sn85_2 78000.000000
Rwneg85_3 in85_3 sn85_3 78000.000000
Rwneg85_4 in85_4 sn85_4 202000.000000
Rwneg85_5 in85_5 sn85_5 202000.000000
Rwneg85_6 in85_6 sn85_6 202000.000000
Rwneg85_7 in85_7 sn85_7 78000.000000
Rwneg85_8 in85_8 sn85_8 202000.000000
Rwneg85_9 in85_9 sn85_9 78000.000000
Rwneg85_10 in85_10 sn85_10 202000.000000
Rwneg85_11 in85_11 sn85_11 202000.000000
Rwneg85_12 in85_12 sn85_12 202000.000000
Rwneg85_13 in85_13 sn85_13 202000.000000
Rwneg85_14 in85_14 sn85_14 78000.000000
Rwneg85_15 in85_15 sn85_15 202000.000000
Rwneg85_16 in85_16 sn85_16 78000.000000
Rwneg85_17 in85_17 sn85_17 78000.000000
Rwneg85_18 in85_18 sn85_18 202000.000000
Rwneg85_19 in85_19 sn85_19 202000.000000
Rwneg85_20 in85_20 sn85_20 202000.000000
Rwneg85_21 in85_21 sn85_21 202000.000000
Rwneg85_22 in85_22 sn85_22 202000.000000
Rwneg85_23 in85_23 sn85_23 202000.000000
Rwneg85_24 in85_24 sn85_24 78000.000000
Rwneg85_25 in85_25 sn85_25 202000.000000
Rwneg85_26 in85_26 sn85_26 202000.000000
Rwneg85_27 in85_27 sn85_27 202000.000000
Rwneg85_28 in85_28 sn85_28 202000.000000
Rwneg85_29 in85_29 sn85_29 78000.000000
Rwneg85_30 in85_30 sn85_30 78000.000000
Rwneg85_31 in85_31 sn85_31 202000.000000
Rwneg85_32 in85_32 sn85_32 78000.000000
Rwneg85_33 in85_33 sn85_33 78000.000000
Rwneg85_34 in85_34 sn85_34 202000.000000
Rwneg85_35 in85_35 sn85_35 202000.000000
Rwneg85_36 in85_36 sn85_36 202000.000000
Rwneg85_37 in85_37 sn85_37 78000.000000
Rwneg85_38 in85_38 sn85_38 202000.000000
Rwneg85_39 in85_39 sn85_39 202000.000000
Rwneg85_40 in85_40 sn85_40 202000.000000
Rwneg85_41 in85_41 sn85_41 78000.000000
Rwneg85_42 in85_42 sn85_42 78000.000000
Rwneg85_43 in85_43 sn85_43 202000.000000
Rwneg85_44 in85_44 sn85_44 78000.000000
Rwneg85_45 in85_45 sn85_45 202000.000000
Rwneg85_46 in85_46 sn85_46 78000.000000
Rwneg85_47 in85_47 sn85_47 202000.000000
Rwneg85_48 in85_48 sn85_48 78000.000000
Rwneg85_49 in85_49 sn85_49 78000.000000
Rwneg85_50 in85_50 sn85_50 202000.000000
Rwneg85_51 in85_51 sn85_51 202000.000000
Rwneg85_52 in85_52 sn85_52 78000.000000
Rwneg85_53 in85_53 sn85_53 202000.000000
Rwneg85_54 in85_54 sn85_54 202000.000000
Rwneg85_55 in85_55 sn85_55 78000.000000
Rwneg85_56 in85_56 sn85_56 202000.000000
Rwneg85_57 in85_57 sn85_57 78000.000000
Rwneg85_58 in85_58 sn85_58 202000.000000
Rwneg85_59 in85_59 sn85_59 78000.000000
Rwneg85_60 in85_60 sn85_60 78000.000000
Rwneg85_61 in85_61 sn85_61 78000.000000
Rwneg85_62 in85_62 sn85_62 202000.000000
Rwneg85_63 in85_63 sn85_63 202000.000000
Rwneg85_64 in85_64 sn85_64 78000.000000
Rwneg85_65 in85_65 sn85_65 78000.000000
Rwneg85_66 in85_66 sn85_66 78000.000000
Rwneg85_67 in85_67 sn85_67 78000.000000
Rwneg85_68 in85_68 sn85_68 78000.000000
Rwneg85_69 in85_69 sn85_69 202000.000000
Rwneg85_70 in85_70 sn85_70 202000.000000
Rwneg85_71 in85_71 sn85_71 202000.000000
Rwneg85_72 in85_72 sn85_72 202000.000000
Rwneg85_73 in85_73 sn85_73 78000.000000
Rwneg85_74 in85_74 sn85_74 78000.000000
Rwneg85_75 in85_75 sn85_75 202000.000000
Rwneg85_76 in85_76 sn85_76 78000.000000
Rwneg85_77 in85_77 sn85_77 202000.000000
Rwneg85_78 in85_78 sn85_78 202000.000000
Rwneg85_79 in85_79 sn85_79 202000.000000
Rwneg85_80 in85_80 sn85_80 202000.000000
Rwneg85_81 in85_81 sn85_81 78000.000000
Rwneg85_82 in85_82 sn85_82 202000.000000
Rwneg85_83 in85_83 sn85_83 78000.000000
Rwneg85_84 in85_84 sn85_84 202000.000000
Rwneg86_1 in86_1 sn86_1 78000.000000
Rwneg86_2 in86_2 sn86_2 202000.000000
Rwneg86_3 in86_3 sn86_3 78000.000000
Rwneg86_4 in86_4 sn86_4 78000.000000
Rwneg86_5 in86_5 sn86_5 78000.000000
Rwneg86_6 in86_6 sn86_6 202000.000000
Rwneg86_7 in86_7 sn86_7 202000.000000
Rwneg86_8 in86_8 sn86_8 78000.000000
Rwneg86_9 in86_9 sn86_9 78000.000000
Rwneg86_10 in86_10 sn86_10 202000.000000
Rwneg86_11 in86_11 sn86_11 78000.000000
Rwneg86_12 in86_12 sn86_12 202000.000000
Rwneg86_13 in86_13 sn86_13 202000.000000
Rwneg86_14 in86_14 sn86_14 202000.000000
Rwneg86_15 in86_15 sn86_15 202000.000000
Rwneg86_16 in86_16 sn86_16 202000.000000
Rwneg86_17 in86_17 sn86_17 202000.000000
Rwneg86_18 in86_18 sn86_18 78000.000000
Rwneg86_19 in86_19 sn86_19 202000.000000
Rwneg86_20 in86_20 sn86_20 78000.000000
Rwneg86_21 in86_21 sn86_21 78000.000000
Rwneg86_22 in86_22 sn86_22 78000.000000
Rwneg86_23 in86_23 sn86_23 78000.000000
Rwneg86_24 in86_24 sn86_24 78000.000000
Rwneg86_25 in86_25 sn86_25 202000.000000
Rwneg86_26 in86_26 sn86_26 78000.000000
Rwneg86_27 in86_27 sn86_27 78000.000000
Rwneg86_28 in86_28 sn86_28 202000.000000
Rwneg86_29 in86_29 sn86_29 78000.000000
Rwneg86_30 in86_30 sn86_30 202000.000000
Rwneg86_31 in86_31 sn86_31 78000.000000
Rwneg86_32 in86_32 sn86_32 202000.000000
Rwneg86_33 in86_33 sn86_33 78000.000000
Rwneg86_34 in86_34 sn86_34 202000.000000
Rwneg86_35 in86_35 sn86_35 78000.000000
Rwneg86_36 in86_36 sn86_36 202000.000000
Rwneg86_37 in86_37 sn86_37 202000.000000
Rwneg86_38 in86_38 sn86_38 202000.000000
Rwneg86_39 in86_39 sn86_39 78000.000000
Rwneg86_40 in86_40 sn86_40 202000.000000
Rwneg86_41 in86_41 sn86_41 78000.000000
Rwneg86_42 in86_42 sn86_42 78000.000000
Rwneg86_43 in86_43 sn86_43 78000.000000
Rwneg86_44 in86_44 sn86_44 202000.000000
Rwneg86_45 in86_45 sn86_45 78000.000000
Rwneg86_46 in86_46 sn86_46 202000.000000
Rwneg86_47 in86_47 sn86_47 202000.000000
Rwneg86_48 in86_48 sn86_48 78000.000000
Rwneg86_49 in86_49 sn86_49 202000.000000
Rwneg86_50 in86_50 sn86_50 202000.000000
Rwneg86_51 in86_51 sn86_51 78000.000000
Rwneg86_52 in86_52 sn86_52 202000.000000
Rwneg86_53 in86_53 sn86_53 78000.000000
Rwneg86_54 in86_54 sn86_54 202000.000000
Rwneg86_55 in86_55 sn86_55 202000.000000
Rwneg86_56 in86_56 sn86_56 78000.000000
Rwneg86_57 in86_57 sn86_57 78000.000000
Rwneg86_58 in86_58 sn86_58 202000.000000
Rwneg86_59 in86_59 sn86_59 78000.000000
Rwneg86_60 in86_60 sn86_60 202000.000000
Rwneg86_61 in86_61 sn86_61 78000.000000
Rwneg86_62 in86_62 sn86_62 78000.000000
Rwneg86_63 in86_63 sn86_63 202000.000000
Rwneg86_64 in86_64 sn86_64 78000.000000
Rwneg86_65 in86_65 sn86_65 78000.000000
Rwneg86_66 in86_66 sn86_66 202000.000000
Rwneg86_67 in86_67 sn86_67 202000.000000
Rwneg86_68 in86_68 sn86_68 202000.000000
Rwneg86_69 in86_69 sn86_69 78000.000000
Rwneg86_70 in86_70 sn86_70 202000.000000
Rwneg86_71 in86_71 sn86_71 78000.000000
Rwneg86_72 in86_72 sn86_72 78000.000000
Rwneg86_73 in86_73 sn86_73 202000.000000
Rwneg86_74 in86_74 sn86_74 202000.000000
Rwneg86_75 in86_75 sn86_75 78000.000000
Rwneg86_76 in86_76 sn86_76 202000.000000
Rwneg86_77 in86_77 sn86_77 78000.000000
Rwneg86_78 in86_78 sn86_78 202000.000000
Rwneg86_79 in86_79 sn86_79 202000.000000
Rwneg86_80 in86_80 sn86_80 78000.000000
Rwneg86_81 in86_81 sn86_81 78000.000000
Rwneg86_82 in86_82 sn86_82 78000.000000
Rwneg86_83 in86_83 sn86_83 78000.000000
Rwneg86_84 in86_84 sn86_84 78000.000000
Rwneg87_1 in87_1 sn87_1 78000.000000
Rwneg87_2 in87_2 sn87_2 78000.000000
Rwneg87_3 in87_3 sn87_3 78000.000000
Rwneg87_4 in87_4 sn87_4 202000.000000
Rwneg87_5 in87_5 sn87_5 202000.000000
Rwneg87_6 in87_6 sn87_6 78000.000000
Rwneg87_7 in87_7 sn87_7 202000.000000
Rwneg87_8 in87_8 sn87_8 78000.000000
Rwneg87_9 in87_9 sn87_9 202000.000000
Rwneg87_10 in87_10 sn87_10 78000.000000
Rwneg87_11 in87_11 sn87_11 202000.000000
Rwneg87_12 in87_12 sn87_12 78000.000000
Rwneg87_13 in87_13 sn87_13 202000.000000
Rwneg87_14 in87_14 sn87_14 202000.000000
Rwneg87_15 in87_15 sn87_15 202000.000000
Rwneg87_16 in87_16 sn87_16 202000.000000
Rwneg87_17 in87_17 sn87_17 78000.000000
Rwneg87_18 in87_18 sn87_18 78000.000000
Rwneg87_19 in87_19 sn87_19 78000.000000
Rwneg87_20 in87_20 sn87_20 78000.000000
Rwneg87_21 in87_21 sn87_21 202000.000000
Rwneg87_22 in87_22 sn87_22 78000.000000
Rwneg87_23 in87_23 sn87_23 78000.000000
Rwneg87_24 in87_24 sn87_24 202000.000000
Rwneg87_25 in87_25 sn87_25 202000.000000
Rwneg87_26 in87_26 sn87_26 78000.000000
Rwneg87_27 in87_27 sn87_27 202000.000000
Rwneg87_28 in87_28 sn87_28 202000.000000
Rwneg87_29 in87_29 sn87_29 78000.000000
Rwneg87_30 in87_30 sn87_30 78000.000000
Rwneg87_31 in87_31 sn87_31 78000.000000
Rwneg87_32 in87_32 sn87_32 78000.000000
Rwneg87_33 in87_33 sn87_33 202000.000000
Rwneg87_34 in87_34 sn87_34 78000.000000
Rwneg87_35 in87_35 sn87_35 202000.000000
Rwneg87_36 in87_36 sn87_36 202000.000000
Rwneg87_37 in87_37 sn87_37 202000.000000
Rwneg87_38 in87_38 sn87_38 78000.000000
Rwneg87_39 in87_39 sn87_39 78000.000000
Rwneg87_40 in87_40 sn87_40 78000.000000
Rwneg87_41 in87_41 sn87_41 202000.000000
Rwneg87_42 in87_42 sn87_42 78000.000000
Rwneg87_43 in87_43 sn87_43 78000.000000
Rwneg87_44 in87_44 sn87_44 78000.000000
Rwneg87_45 in87_45 sn87_45 78000.000000
Rwneg87_46 in87_46 sn87_46 202000.000000
Rwneg87_47 in87_47 sn87_47 202000.000000
Rwneg87_48 in87_48 sn87_48 202000.000000
Rwneg87_49 in87_49 sn87_49 202000.000000
Rwneg87_50 in87_50 sn87_50 202000.000000
Rwneg87_51 in87_51 sn87_51 202000.000000
Rwneg87_52 in87_52 sn87_52 202000.000000
Rwneg87_53 in87_53 sn87_53 78000.000000
Rwneg87_54 in87_54 sn87_54 202000.000000
Rwneg87_55 in87_55 sn87_55 78000.000000
Rwneg87_56 in87_56 sn87_56 78000.000000
Rwneg87_57 in87_57 sn87_57 202000.000000
Rwneg87_58 in87_58 sn87_58 78000.000000
Rwneg87_59 in87_59 sn87_59 202000.000000
Rwneg87_60 in87_60 sn87_60 78000.000000
Rwneg87_61 in87_61 sn87_61 78000.000000
Rwneg87_62 in87_62 sn87_62 202000.000000
Rwneg87_63 in87_63 sn87_63 78000.000000
Rwneg87_64 in87_64 sn87_64 78000.000000
Rwneg87_65 in87_65 sn87_65 202000.000000
Rwneg87_66 in87_66 sn87_66 202000.000000
Rwneg87_67 in87_67 sn87_67 202000.000000
Rwneg87_68 in87_68 sn87_68 78000.000000
Rwneg87_69 in87_69 sn87_69 78000.000000
Rwneg87_70 in87_70 sn87_70 202000.000000
Rwneg87_71 in87_71 sn87_71 78000.000000
Rwneg87_72 in87_72 sn87_72 78000.000000
Rwneg87_73 in87_73 sn87_73 78000.000000
Rwneg87_74 in87_74 sn87_74 78000.000000
Rwneg87_75 in87_75 sn87_75 202000.000000
Rwneg87_76 in87_76 sn87_76 202000.000000
Rwneg87_77 in87_77 sn87_77 78000.000000
Rwneg87_78 in87_78 sn87_78 202000.000000
Rwneg87_79 in87_79 sn87_79 78000.000000
Rwneg87_80 in87_80 sn87_80 202000.000000
Rwneg87_81 in87_81 sn87_81 78000.000000
Rwneg87_82 in87_82 sn87_82 202000.000000
Rwneg87_83 in87_83 sn87_83 78000.000000
Rwneg87_84 in87_84 sn87_84 78000.000000
Rwneg88_1 in88_1 sn88_1 78000.000000
Rwneg88_2 in88_2 sn88_2 202000.000000
Rwneg88_3 in88_3 sn88_3 202000.000000
Rwneg88_4 in88_4 sn88_4 78000.000000
Rwneg88_5 in88_5 sn88_5 202000.000000
Rwneg88_6 in88_6 sn88_6 202000.000000
Rwneg88_7 in88_7 sn88_7 202000.000000
Rwneg88_8 in88_8 sn88_8 78000.000000
Rwneg88_9 in88_9 sn88_9 78000.000000
Rwneg88_10 in88_10 sn88_10 78000.000000
Rwneg88_11 in88_11 sn88_11 202000.000000
Rwneg88_12 in88_12 sn88_12 78000.000000
Rwneg88_13 in88_13 sn88_13 78000.000000
Rwneg88_14 in88_14 sn88_14 202000.000000
Rwneg88_15 in88_15 sn88_15 202000.000000
Rwneg88_16 in88_16 sn88_16 202000.000000
Rwneg88_17 in88_17 sn88_17 202000.000000
Rwneg88_18 in88_18 sn88_18 78000.000000
Rwneg88_19 in88_19 sn88_19 202000.000000
Rwneg88_20 in88_20 sn88_20 78000.000000
Rwneg88_21 in88_21 sn88_21 78000.000000
Rwneg88_22 in88_22 sn88_22 202000.000000
Rwneg88_23 in88_23 sn88_23 202000.000000
Rwneg88_24 in88_24 sn88_24 202000.000000
Rwneg88_25 in88_25 sn88_25 202000.000000
Rwneg88_26 in88_26 sn88_26 78000.000000
Rwneg88_27 in88_27 sn88_27 202000.000000
Rwneg88_28 in88_28 sn88_28 78000.000000
Rwneg88_29 in88_29 sn88_29 78000.000000
Rwneg88_30 in88_30 sn88_30 78000.000000
Rwneg88_31 in88_31 sn88_31 78000.000000
Rwneg88_32 in88_32 sn88_32 202000.000000
Rwneg88_33 in88_33 sn88_33 202000.000000
Rwneg88_34 in88_34 sn88_34 78000.000000
Rwneg88_35 in88_35 sn88_35 78000.000000
Rwneg88_36 in88_36 sn88_36 202000.000000
Rwneg88_37 in88_37 sn88_37 78000.000000
Rwneg88_38 in88_38 sn88_38 202000.000000
Rwneg88_39 in88_39 sn88_39 78000.000000
Rwneg88_40 in88_40 sn88_40 202000.000000
Rwneg88_41 in88_41 sn88_41 78000.000000
Rwneg88_42 in88_42 sn88_42 202000.000000
Rwneg88_43 in88_43 sn88_43 78000.000000
Rwneg88_44 in88_44 sn88_44 202000.000000
Rwneg88_45 in88_45 sn88_45 78000.000000
Rwneg88_46 in88_46 sn88_46 202000.000000
Rwneg88_47 in88_47 sn88_47 202000.000000
Rwneg88_48 in88_48 sn88_48 78000.000000
Rwneg88_49 in88_49 sn88_49 78000.000000
Rwneg88_50 in88_50 sn88_50 78000.000000
Rwneg88_51 in88_51 sn88_51 78000.000000
Rwneg88_52 in88_52 sn88_52 78000.000000
Rwneg88_53 in88_53 sn88_53 202000.000000
Rwneg88_54 in88_54 sn88_54 78000.000000
Rwneg88_55 in88_55 sn88_55 202000.000000
Rwneg88_56 in88_56 sn88_56 78000.000000
Rwneg88_57 in88_57 sn88_57 78000.000000
Rwneg88_58 in88_58 sn88_58 202000.000000
Rwneg88_59 in88_59 sn88_59 78000.000000
Rwneg88_60 in88_60 sn88_60 202000.000000
Rwneg88_61 in88_61 sn88_61 78000.000000
Rwneg88_62 in88_62 sn88_62 202000.000000
Rwneg88_63 in88_63 sn88_63 78000.000000
Rwneg88_64 in88_64 sn88_64 78000.000000
Rwneg88_65 in88_65 sn88_65 78000.000000
Rwneg88_66 in88_66 sn88_66 78000.000000
Rwneg88_67 in88_67 sn88_67 202000.000000
Rwneg88_68 in88_68 sn88_68 202000.000000
Rwneg88_69 in88_69 sn88_69 78000.000000
Rwneg88_70 in88_70 sn88_70 78000.000000
Rwneg88_71 in88_71 sn88_71 78000.000000
Rwneg88_72 in88_72 sn88_72 202000.000000
Rwneg88_73 in88_73 sn88_73 78000.000000
Rwneg88_74 in88_74 sn88_74 202000.000000
Rwneg88_75 in88_75 sn88_75 78000.000000
Rwneg88_76 in88_76 sn88_76 78000.000000
Rwneg88_77 in88_77 sn88_77 78000.000000
Rwneg88_78 in88_78 sn88_78 202000.000000
Rwneg88_79 in88_79 sn88_79 78000.000000
Rwneg88_80 in88_80 sn88_80 78000.000000
Rwneg88_81 in88_81 sn88_81 202000.000000
Rwneg88_82 in88_82 sn88_82 78000.000000
Rwneg88_83 in88_83 sn88_83 202000.000000
Rwneg88_84 in88_84 sn88_84 78000.000000
Rwneg89_1 in89_1 sn89_1 78000.000000
Rwneg89_2 in89_2 sn89_2 78000.000000
Rwneg89_3 in89_3 sn89_3 78000.000000
Rwneg89_4 in89_4 sn89_4 78000.000000
Rwneg89_5 in89_5 sn89_5 202000.000000
Rwneg89_6 in89_6 sn89_6 78000.000000
Rwneg89_7 in89_7 sn89_7 202000.000000
Rwneg89_8 in89_8 sn89_8 78000.000000
Rwneg89_9 in89_9 sn89_9 78000.000000
Rwneg89_10 in89_10 sn89_10 202000.000000
Rwneg89_11 in89_11 sn89_11 78000.000000
Rwneg89_12 in89_12 sn89_12 78000.000000
Rwneg89_13 in89_13 sn89_13 202000.000000
Rwneg89_14 in89_14 sn89_14 202000.000000
Rwneg89_15 in89_15 sn89_15 202000.000000
Rwneg89_16 in89_16 sn89_16 78000.000000
Rwneg89_17 in89_17 sn89_17 202000.000000
Rwneg89_18 in89_18 sn89_18 78000.000000
Rwneg89_19 in89_19 sn89_19 78000.000000
Rwneg89_20 in89_20 sn89_20 78000.000000
Rwneg89_21 in89_21 sn89_21 78000.000000
Rwneg89_22 in89_22 sn89_22 202000.000000
Rwneg89_23 in89_23 sn89_23 202000.000000
Rwneg89_24 in89_24 sn89_24 202000.000000
Rwneg89_25 in89_25 sn89_25 202000.000000
Rwneg89_26 in89_26 sn89_26 78000.000000
Rwneg89_27 in89_27 sn89_27 202000.000000
Rwneg89_28 in89_28 sn89_28 78000.000000
Rwneg89_29 in89_29 sn89_29 202000.000000
Rwneg89_30 in89_30 sn89_30 202000.000000
Rwneg89_31 in89_31 sn89_31 202000.000000
Rwneg89_32 in89_32 sn89_32 78000.000000
Rwneg89_33 in89_33 sn89_33 202000.000000
Rwneg89_34 in89_34 sn89_34 78000.000000
Rwneg89_35 in89_35 sn89_35 202000.000000
Rwneg89_36 in89_36 sn89_36 78000.000000
Rwneg89_37 in89_37 sn89_37 78000.000000
Rwneg89_38 in89_38 sn89_38 78000.000000
Rwneg89_39 in89_39 sn89_39 78000.000000
Rwneg89_40 in89_40 sn89_40 202000.000000
Rwneg89_41 in89_41 sn89_41 78000.000000
Rwneg89_42 in89_42 sn89_42 78000.000000
Rwneg89_43 in89_43 sn89_43 202000.000000
Rwneg89_44 in89_44 sn89_44 78000.000000
Rwneg89_45 in89_45 sn89_45 78000.000000
Rwneg89_46 in89_46 sn89_46 202000.000000
Rwneg89_47 in89_47 sn89_47 78000.000000
Rwneg89_48 in89_48 sn89_48 78000.000000
Rwneg89_49 in89_49 sn89_49 78000.000000
Rwneg89_50 in89_50 sn89_50 78000.000000
Rwneg89_51 in89_51 sn89_51 202000.000000
Rwneg89_52 in89_52 sn89_52 78000.000000
Rwneg89_53 in89_53 sn89_53 202000.000000
Rwneg89_54 in89_54 sn89_54 202000.000000
Rwneg89_55 in89_55 sn89_55 78000.000000
Rwneg89_56 in89_56 sn89_56 78000.000000
Rwneg89_57 in89_57 sn89_57 202000.000000
Rwneg89_58 in89_58 sn89_58 202000.000000
Rwneg89_59 in89_59 sn89_59 202000.000000
Rwneg89_60 in89_60 sn89_60 202000.000000
Rwneg89_61 in89_61 sn89_61 78000.000000
Rwneg89_62 in89_62 sn89_62 202000.000000
Rwneg89_63 in89_63 sn89_63 78000.000000
Rwneg89_64 in89_64 sn89_64 78000.000000
Rwneg89_65 in89_65 sn89_65 78000.000000
Rwneg89_66 in89_66 sn89_66 202000.000000
Rwneg89_67 in89_67 sn89_67 202000.000000
Rwneg89_68 in89_68 sn89_68 202000.000000
Rwneg89_69 in89_69 sn89_69 78000.000000
Rwneg89_70 in89_70 sn89_70 202000.000000
Rwneg89_71 in89_71 sn89_71 78000.000000
Rwneg89_72 in89_72 sn89_72 202000.000000
Rwneg89_73 in89_73 sn89_73 202000.000000
Rwneg89_74 in89_74 sn89_74 202000.000000
Rwneg89_75 in89_75 sn89_75 78000.000000
Rwneg89_76 in89_76 sn89_76 78000.000000
Rwneg89_77 in89_77 sn89_77 78000.000000
Rwneg89_78 in89_78 sn89_78 78000.000000
Rwneg89_79 in89_79 sn89_79 78000.000000
Rwneg89_80 in89_80 sn89_80 202000.000000
Rwneg89_81 in89_81 sn89_81 202000.000000
Rwneg89_82 in89_82 sn89_82 78000.000000
Rwneg89_83 in89_83 sn89_83 202000.000000
Rwneg89_84 in89_84 sn89_84 78000.000000
Rwneg90_1 in90_1 sn90_1 78000.000000
Rwneg90_2 in90_2 sn90_2 202000.000000
Rwneg90_3 in90_3 sn90_3 202000.000000
Rwneg90_4 in90_4 sn90_4 202000.000000
Rwneg90_5 in90_5 sn90_5 78000.000000
Rwneg90_6 in90_6 sn90_6 202000.000000
Rwneg90_7 in90_7 sn90_7 78000.000000
Rwneg90_8 in90_8 sn90_8 202000.000000
Rwneg90_9 in90_9 sn90_9 78000.000000
Rwneg90_10 in90_10 sn90_10 202000.000000
Rwneg90_11 in90_11 sn90_11 78000.000000
Rwneg90_12 in90_12 sn90_12 202000.000000
Rwneg90_13 in90_13 sn90_13 202000.000000
Rwneg90_14 in90_14 sn90_14 202000.000000
Rwneg90_15 in90_15 sn90_15 202000.000000
Rwneg90_16 in90_16 sn90_16 78000.000000
Rwneg90_17 in90_17 sn90_17 202000.000000
Rwneg90_18 in90_18 sn90_18 78000.000000
Rwneg90_19 in90_19 sn90_19 78000.000000
Rwneg90_20 in90_20 sn90_20 78000.000000
Rwneg90_21 in90_21 sn90_21 202000.000000
Rwneg90_22 in90_22 sn90_22 202000.000000
Rwneg90_23 in90_23 sn90_23 202000.000000
Rwneg90_24 in90_24 sn90_24 202000.000000
Rwneg90_25 in90_25 sn90_25 202000.000000
Rwneg90_26 in90_26 sn90_26 202000.000000
Rwneg90_27 in90_27 sn90_27 202000.000000
Rwneg90_28 in90_28 sn90_28 78000.000000
Rwneg90_29 in90_29 sn90_29 78000.000000
Rwneg90_30 in90_30 sn90_30 78000.000000
Rwneg90_31 in90_31 sn90_31 202000.000000
Rwneg90_32 in90_32 sn90_32 78000.000000
Rwneg90_33 in90_33 sn90_33 78000.000000
Rwneg90_34 in90_34 sn90_34 78000.000000
Rwneg90_35 in90_35 sn90_35 202000.000000
Rwneg90_36 in90_36 sn90_36 202000.000000
Rwneg90_37 in90_37 sn90_37 78000.000000
Rwneg90_38 in90_38 sn90_38 78000.000000
Rwneg90_39 in90_39 sn90_39 78000.000000
Rwneg90_40 in90_40 sn90_40 78000.000000
Rwneg90_41 in90_41 sn90_41 202000.000000
Rwneg90_42 in90_42 sn90_42 78000.000000
Rwneg90_43 in90_43 sn90_43 202000.000000
Rwneg90_44 in90_44 sn90_44 202000.000000
Rwneg90_45 in90_45 sn90_45 78000.000000
Rwneg90_46 in90_46 sn90_46 202000.000000
Rwneg90_47 in90_47 sn90_47 202000.000000
Rwneg90_48 in90_48 sn90_48 78000.000000
Rwneg90_49 in90_49 sn90_49 78000.000000
Rwneg90_50 in90_50 sn90_50 78000.000000
Rwneg90_51 in90_51 sn90_51 202000.000000
Rwneg90_52 in90_52 sn90_52 78000.000000
Rwneg90_53 in90_53 sn90_53 78000.000000
Rwneg90_54 in90_54 sn90_54 202000.000000
Rwneg90_55 in90_55 sn90_55 78000.000000
Rwneg90_56 in90_56 sn90_56 78000.000000
Rwneg90_57 in90_57 sn90_57 78000.000000
Rwneg90_58 in90_58 sn90_58 202000.000000
Rwneg90_59 in90_59 sn90_59 202000.000000
Rwneg90_60 in90_60 sn90_60 202000.000000
Rwneg90_61 in90_61 sn90_61 202000.000000
Rwneg90_62 in90_62 sn90_62 202000.000000
Rwneg90_63 in90_63 sn90_63 202000.000000
Rwneg90_64 in90_64 sn90_64 78000.000000
Rwneg90_65 in90_65 sn90_65 202000.000000
Rwneg90_66 in90_66 sn90_66 78000.000000
Rwneg90_67 in90_67 sn90_67 202000.000000
Rwneg90_68 in90_68 sn90_68 202000.000000
Rwneg90_69 in90_69 sn90_69 78000.000000
Rwneg90_70 in90_70 sn90_70 202000.000000
Rwneg90_71 in90_71 sn90_71 78000.000000
Rwneg90_72 in90_72 sn90_72 202000.000000
Rwneg90_73 in90_73 sn90_73 202000.000000
Rwneg90_74 in90_74 sn90_74 202000.000000
Rwneg90_75 in90_75 sn90_75 78000.000000
Rwneg90_76 in90_76 sn90_76 202000.000000
Rwneg90_77 in90_77 sn90_77 202000.000000
Rwneg90_78 in90_78 sn90_78 202000.000000
Rwneg90_79 in90_79 sn90_79 78000.000000
Rwneg90_80 in90_80 sn90_80 202000.000000
Rwneg90_81 in90_81 sn90_81 202000.000000
Rwneg90_82 in90_82 sn90_82 202000.000000
Rwneg90_83 in90_83 sn90_83 202000.000000
Rwneg90_84 in90_84 sn90_84 202000.000000
Rwneg91_1 in91_1 sn91_1 202000.000000
Rwneg91_2 in91_2 sn91_2 202000.000000
Rwneg91_3 in91_3 sn91_3 78000.000000
Rwneg91_4 in91_4 sn91_4 78000.000000
Rwneg91_5 in91_5 sn91_5 78000.000000
Rwneg91_6 in91_6 sn91_6 202000.000000
Rwneg91_7 in91_7 sn91_7 202000.000000
Rwneg91_8 in91_8 sn91_8 202000.000000
Rwneg91_9 in91_9 sn91_9 202000.000000
Rwneg91_10 in91_10 sn91_10 202000.000000
Rwneg91_11 in91_11 sn91_11 202000.000000
Rwneg91_12 in91_12 sn91_12 202000.000000
Rwneg91_13 in91_13 sn91_13 78000.000000
Rwneg91_14 in91_14 sn91_14 78000.000000
Rwneg91_15 in91_15 sn91_15 202000.000000
Rwneg91_16 in91_16 sn91_16 202000.000000
Rwneg91_17 in91_17 sn91_17 202000.000000
Rwneg91_18 in91_18 sn91_18 202000.000000
Rwneg91_19 in91_19 sn91_19 202000.000000
Rwneg91_20 in91_20 sn91_20 78000.000000
Rwneg91_21 in91_21 sn91_21 202000.000000
Rwneg91_22 in91_22 sn91_22 202000.000000
Rwneg91_23 in91_23 sn91_23 78000.000000
Rwneg91_24 in91_24 sn91_24 202000.000000
Rwneg91_25 in91_25 sn91_25 202000.000000
Rwneg91_26 in91_26 sn91_26 78000.000000
Rwneg91_27 in91_27 sn91_27 202000.000000
Rwneg91_28 in91_28 sn91_28 202000.000000
Rwneg91_29 in91_29 sn91_29 78000.000000
Rwneg91_30 in91_30 sn91_30 202000.000000
Rwneg91_31 in91_31 sn91_31 78000.000000
Rwneg91_32 in91_32 sn91_32 202000.000000
Rwneg91_33 in91_33 sn91_33 202000.000000
Rwneg91_34 in91_34 sn91_34 78000.000000
Rwneg91_35 in91_35 sn91_35 78000.000000
Rwneg91_36 in91_36 sn91_36 78000.000000
Rwneg91_37 in91_37 sn91_37 202000.000000
Rwneg91_38 in91_38 sn91_38 78000.000000
Rwneg91_39 in91_39 sn91_39 78000.000000
Rwneg91_40 in91_40 sn91_40 202000.000000
Rwneg91_41 in91_41 sn91_41 202000.000000
Rwneg91_42 in91_42 sn91_42 78000.000000
Rwneg91_43 in91_43 sn91_43 202000.000000
Rwneg91_44 in91_44 sn91_44 202000.000000
Rwneg91_45 in91_45 sn91_45 202000.000000
Rwneg91_46 in91_46 sn91_46 78000.000000
Rwneg91_47 in91_47 sn91_47 78000.000000
Rwneg91_48 in91_48 sn91_48 78000.000000
Rwneg91_49 in91_49 sn91_49 78000.000000
Rwneg91_50 in91_50 sn91_50 78000.000000
Rwneg91_51 in91_51 sn91_51 78000.000000
Rwneg91_52 in91_52 sn91_52 78000.000000
Rwneg91_53 in91_53 sn91_53 78000.000000
Rwneg91_54 in91_54 sn91_54 202000.000000
Rwneg91_55 in91_55 sn91_55 202000.000000
Rwneg91_56 in91_56 sn91_56 202000.000000
Rwneg91_57 in91_57 sn91_57 78000.000000
Rwneg91_58 in91_58 sn91_58 202000.000000
Rwneg91_59 in91_59 sn91_59 78000.000000
Rwneg91_60 in91_60 sn91_60 78000.000000
Rwneg91_61 in91_61 sn91_61 202000.000000
Rwneg91_62 in91_62 sn91_62 202000.000000
Rwneg91_63 in91_63 sn91_63 202000.000000
Rwneg91_64 in91_64 sn91_64 78000.000000
Rwneg91_65 in91_65 sn91_65 202000.000000
Rwneg91_66 in91_66 sn91_66 202000.000000
Rwneg91_67 in91_67 sn91_67 78000.000000
Rwneg91_68 in91_68 sn91_68 202000.000000
Rwneg91_69 in91_69 sn91_69 202000.000000
Rwneg91_70 in91_70 sn91_70 78000.000000
Rwneg91_71 in91_71 sn91_71 202000.000000
Rwneg91_72 in91_72 sn91_72 202000.000000
Rwneg91_73 in91_73 sn91_73 202000.000000
Rwneg91_74 in91_74 sn91_74 78000.000000
Rwneg91_75 in91_75 sn91_75 78000.000000
Rwneg91_76 in91_76 sn91_76 78000.000000
Rwneg91_77 in91_77 sn91_77 202000.000000
Rwneg91_78 in91_78 sn91_78 78000.000000
Rwneg91_79 in91_79 sn91_79 78000.000000
Rwneg91_80 in91_80 sn91_80 202000.000000
Rwneg91_81 in91_81 sn91_81 78000.000000
Rwneg91_82 in91_82 sn91_82 202000.000000
Rwneg91_83 in91_83 sn91_83 78000.000000
Rwneg91_84 in91_84 sn91_84 78000.000000
Rwneg92_1 in92_1 sn92_1 78000.000000
Rwneg92_2 in92_2 sn92_2 202000.000000
Rwneg92_3 in92_3 sn92_3 202000.000000
Rwneg92_4 in92_4 sn92_4 78000.000000
Rwneg92_5 in92_5 sn92_5 78000.000000
Rwneg92_6 in92_6 sn92_6 202000.000000
Rwneg92_7 in92_7 sn92_7 202000.000000
Rwneg92_8 in92_8 sn92_8 202000.000000
Rwneg92_9 in92_9 sn92_9 78000.000000
Rwneg92_10 in92_10 sn92_10 78000.000000
Rwneg92_11 in92_11 sn92_11 78000.000000
Rwneg92_12 in92_12 sn92_12 78000.000000
Rwneg92_13 in92_13 sn92_13 78000.000000
Rwneg92_14 in92_14 sn92_14 202000.000000
Rwneg92_15 in92_15 sn92_15 202000.000000
Rwneg92_16 in92_16 sn92_16 78000.000000
Rwneg92_17 in92_17 sn92_17 202000.000000
Rwneg92_18 in92_18 sn92_18 202000.000000
Rwneg92_19 in92_19 sn92_19 78000.000000
Rwneg92_20 in92_20 sn92_20 202000.000000
Rwneg92_21 in92_21 sn92_21 78000.000000
Rwneg92_22 in92_22 sn92_22 78000.000000
Rwneg92_23 in92_23 sn92_23 202000.000000
Rwneg92_24 in92_24 sn92_24 202000.000000
Rwneg92_25 in92_25 sn92_25 202000.000000
Rwneg92_26 in92_26 sn92_26 78000.000000
Rwneg92_27 in92_27 sn92_27 78000.000000
Rwneg92_28 in92_28 sn92_28 202000.000000
Rwneg92_29 in92_29 sn92_29 78000.000000
Rwneg92_30 in92_30 sn92_30 202000.000000
Rwneg92_31 in92_31 sn92_31 78000.000000
Rwneg92_32 in92_32 sn92_32 202000.000000
Rwneg92_33 in92_33 sn92_33 202000.000000
Rwneg92_34 in92_34 sn92_34 78000.000000
Rwneg92_35 in92_35 sn92_35 202000.000000
Rwneg92_36 in92_36 sn92_36 202000.000000
Rwneg92_37 in92_37 sn92_37 78000.000000
Rwneg92_38 in92_38 sn92_38 78000.000000
Rwneg92_39 in92_39 sn92_39 78000.000000
Rwneg92_40 in92_40 sn92_40 78000.000000
Rwneg92_41 in92_41 sn92_41 202000.000000
Rwneg92_42 in92_42 sn92_42 202000.000000
Rwneg92_43 in92_43 sn92_43 78000.000000
Rwneg92_44 in92_44 sn92_44 202000.000000
Rwneg92_45 in92_45 sn92_45 202000.000000
Rwneg92_46 in92_46 sn92_46 202000.000000
Rwneg92_47 in92_47 sn92_47 202000.000000
Rwneg92_48 in92_48 sn92_48 202000.000000
Rwneg92_49 in92_49 sn92_49 78000.000000
Rwneg92_50 in92_50 sn92_50 78000.000000
Rwneg92_51 in92_51 sn92_51 78000.000000
Rwneg92_52 in92_52 sn92_52 78000.000000
Rwneg92_53 in92_53 sn92_53 78000.000000
Rwneg92_54 in92_54 sn92_54 78000.000000
Rwneg92_55 in92_55 sn92_55 202000.000000
Rwneg92_56 in92_56 sn92_56 202000.000000
Rwneg92_57 in92_57 sn92_57 202000.000000
Rwneg92_58 in92_58 sn92_58 202000.000000
Rwneg92_59 in92_59 sn92_59 78000.000000
Rwneg92_60 in92_60 sn92_60 78000.000000
Rwneg92_61 in92_61 sn92_61 202000.000000
Rwneg92_62 in92_62 sn92_62 78000.000000
Rwneg92_63 in92_63 sn92_63 202000.000000
Rwneg92_64 in92_64 sn92_64 78000.000000
Rwneg92_65 in92_65 sn92_65 78000.000000
Rwneg92_66 in92_66 sn92_66 78000.000000
Rwneg92_67 in92_67 sn92_67 78000.000000
Rwneg92_68 in92_68 sn92_68 202000.000000
Rwneg92_69 in92_69 sn92_69 78000.000000
Rwneg92_70 in92_70 sn92_70 202000.000000
Rwneg92_71 in92_71 sn92_71 202000.000000
Rwneg92_72 in92_72 sn92_72 202000.000000
Rwneg92_73 in92_73 sn92_73 78000.000000
Rwneg92_74 in92_74 sn92_74 202000.000000
Rwneg92_75 in92_75 sn92_75 202000.000000
Rwneg92_76 in92_76 sn92_76 202000.000000
Rwneg92_77 in92_77 sn92_77 202000.000000
Rwneg92_78 in92_78 sn92_78 202000.000000
Rwneg92_79 in92_79 sn92_79 202000.000000
Rwneg92_80 in92_80 sn92_80 202000.000000
Rwneg92_81 in92_81 sn92_81 202000.000000
Rwneg92_82 in92_82 sn92_82 202000.000000
Rwneg92_83 in92_83 sn92_83 202000.000000
Rwneg92_84 in92_84 sn92_84 202000.000000
Rwneg93_1 in93_1 sn93_1 202000.000000
Rwneg93_2 in93_2 sn93_2 78000.000000
Rwneg93_3 in93_3 sn93_3 78000.000000
Rwneg93_4 in93_4 sn93_4 78000.000000
Rwneg93_5 in93_5 sn93_5 78000.000000
Rwneg93_6 in93_6 sn93_6 78000.000000
Rwneg93_7 in93_7 sn93_7 202000.000000
Rwneg93_8 in93_8 sn93_8 202000.000000
Rwneg93_9 in93_9 sn93_9 202000.000000
Rwneg93_10 in93_10 sn93_10 202000.000000
Rwneg93_11 in93_11 sn93_11 202000.000000
Rwneg93_12 in93_12 sn93_12 202000.000000
Rwneg93_13 in93_13 sn93_13 202000.000000
Rwneg93_14 in93_14 sn93_14 202000.000000
Rwneg93_15 in93_15 sn93_15 202000.000000
Rwneg93_16 in93_16 sn93_16 202000.000000
Rwneg93_17 in93_17 sn93_17 202000.000000
Rwneg93_18 in93_18 sn93_18 202000.000000
Rwneg93_19 in93_19 sn93_19 78000.000000
Rwneg93_20 in93_20 sn93_20 78000.000000
Rwneg93_21 in93_21 sn93_21 202000.000000
Rwneg93_22 in93_22 sn93_22 78000.000000
Rwneg93_23 in93_23 sn93_23 78000.000000
Rwneg93_24 in93_24 sn93_24 202000.000000
Rwneg93_25 in93_25 sn93_25 78000.000000
Rwneg93_26 in93_26 sn93_26 202000.000000
Rwneg93_27 in93_27 sn93_27 202000.000000
Rwneg93_28 in93_28 sn93_28 202000.000000
Rwneg93_29 in93_29 sn93_29 78000.000000
Rwneg93_30 in93_30 sn93_30 78000.000000
Rwneg93_31 in93_31 sn93_31 202000.000000
Rwneg93_32 in93_32 sn93_32 202000.000000
Rwneg93_33 in93_33 sn93_33 78000.000000
Rwneg93_34 in93_34 sn93_34 202000.000000
Rwneg93_35 in93_35 sn93_35 78000.000000
Rwneg93_36 in93_36 sn93_36 202000.000000
Rwneg93_37 in93_37 sn93_37 202000.000000
Rwneg93_38 in93_38 sn93_38 78000.000000
Rwneg93_39 in93_39 sn93_39 202000.000000
Rwneg93_40 in93_40 sn93_40 78000.000000
Rwneg93_41 in93_41 sn93_41 78000.000000
Rwneg93_42 in93_42 sn93_42 78000.000000
Rwneg93_43 in93_43 sn93_43 202000.000000
Rwneg93_44 in93_44 sn93_44 202000.000000
Rwneg93_45 in93_45 sn93_45 78000.000000
Rwneg93_46 in93_46 sn93_46 202000.000000
Rwneg93_47 in93_47 sn93_47 78000.000000
Rwneg93_48 in93_48 sn93_48 202000.000000
Rwneg93_49 in93_49 sn93_49 78000.000000
Rwneg93_50 in93_50 sn93_50 202000.000000
Rwneg93_51 in93_51 sn93_51 78000.000000
Rwneg93_52 in93_52 sn93_52 202000.000000
Rwneg93_53 in93_53 sn93_53 202000.000000
Rwneg93_54 in93_54 sn93_54 202000.000000
Rwneg93_55 in93_55 sn93_55 202000.000000
Rwneg93_56 in93_56 sn93_56 78000.000000
Rwneg93_57 in93_57 sn93_57 78000.000000
Rwneg93_58 in93_58 sn93_58 78000.000000
Rwneg93_59 in93_59 sn93_59 202000.000000
Rwneg93_60 in93_60 sn93_60 202000.000000
Rwneg93_61 in93_61 sn93_61 202000.000000
Rwneg93_62 in93_62 sn93_62 202000.000000
Rwneg93_63 in93_63 sn93_63 202000.000000
Rwneg93_64 in93_64 sn93_64 202000.000000
Rwneg93_65 in93_65 sn93_65 78000.000000
Rwneg93_66 in93_66 sn93_66 202000.000000
Rwneg93_67 in93_67 sn93_67 202000.000000
Rwneg93_68 in93_68 sn93_68 202000.000000
Rwneg93_69 in93_69 sn93_69 202000.000000
Rwneg93_70 in93_70 sn93_70 78000.000000
Rwneg93_71 in93_71 sn93_71 202000.000000
Rwneg93_72 in93_72 sn93_72 202000.000000
Rwneg93_73 in93_73 sn93_73 202000.000000
Rwneg93_74 in93_74 sn93_74 78000.000000
Rwneg93_75 in93_75 sn93_75 78000.000000
Rwneg93_76 in93_76 sn93_76 202000.000000
Rwneg93_77 in93_77 sn93_77 78000.000000
Rwneg93_78 in93_78 sn93_78 78000.000000
Rwneg93_79 in93_79 sn93_79 202000.000000
Rwneg93_80 in93_80 sn93_80 202000.000000
Rwneg93_81 in93_81 sn93_81 78000.000000
Rwneg93_82 in93_82 sn93_82 202000.000000
Rwneg93_83 in93_83 sn93_83 78000.000000
Rwneg93_84 in93_84 sn93_84 78000.000000
Rwneg94_1 in94_1 sn94_1 78000.000000
Rwneg94_2 in94_2 sn94_2 78000.000000
Rwneg94_3 in94_3 sn94_3 202000.000000
Rwneg94_4 in94_4 sn94_4 202000.000000
Rwneg94_5 in94_5 sn94_5 202000.000000
Rwneg94_6 in94_6 sn94_6 202000.000000
Rwneg94_7 in94_7 sn94_7 78000.000000
Rwneg94_8 in94_8 sn94_8 78000.000000
Rwneg94_9 in94_9 sn94_9 202000.000000
Rwneg94_10 in94_10 sn94_10 202000.000000
Rwneg94_11 in94_11 sn94_11 202000.000000
Rwneg94_12 in94_12 sn94_12 202000.000000
Rwneg94_13 in94_13 sn94_13 78000.000000
Rwneg94_14 in94_14 sn94_14 202000.000000
Rwneg94_15 in94_15 sn94_15 202000.000000
Rwneg94_16 in94_16 sn94_16 78000.000000
Rwneg94_17 in94_17 sn94_17 78000.000000
Rwneg94_18 in94_18 sn94_18 202000.000000
Rwneg94_19 in94_19 sn94_19 202000.000000
Rwneg94_20 in94_20 sn94_20 78000.000000
Rwneg94_21 in94_21 sn94_21 202000.000000
Rwneg94_22 in94_22 sn94_22 78000.000000
Rwneg94_23 in94_23 sn94_23 78000.000000
Rwneg94_24 in94_24 sn94_24 202000.000000
Rwneg94_25 in94_25 sn94_25 78000.000000
Rwneg94_26 in94_26 sn94_26 202000.000000
Rwneg94_27 in94_27 sn94_27 78000.000000
Rwneg94_28 in94_28 sn94_28 78000.000000
Rwneg94_29 in94_29 sn94_29 202000.000000
Rwneg94_30 in94_30 sn94_30 202000.000000
Rwneg94_31 in94_31 sn94_31 202000.000000
Rwneg94_32 in94_32 sn94_32 202000.000000
Rwneg94_33 in94_33 sn94_33 78000.000000
Rwneg94_34 in94_34 sn94_34 202000.000000
Rwneg94_35 in94_35 sn94_35 78000.000000
Rwneg94_36 in94_36 sn94_36 202000.000000
Rwneg94_37 in94_37 sn94_37 202000.000000
Rwneg94_38 in94_38 sn94_38 202000.000000
Rwneg94_39 in94_39 sn94_39 202000.000000
Rwneg94_40 in94_40 sn94_40 78000.000000
Rwneg94_41 in94_41 sn94_41 78000.000000
Rwneg94_42 in94_42 sn94_42 78000.000000
Rwneg94_43 in94_43 sn94_43 202000.000000
Rwneg94_44 in94_44 sn94_44 78000.000000
Rwneg94_45 in94_45 sn94_45 78000.000000
Rwneg94_46 in94_46 sn94_46 202000.000000
Rwneg94_47 in94_47 sn94_47 202000.000000
Rwneg94_48 in94_48 sn94_48 78000.000000
Rwneg94_49 in94_49 sn94_49 78000.000000
Rwneg94_50 in94_50 sn94_50 78000.000000
Rwneg94_51 in94_51 sn94_51 78000.000000
Rwneg94_52 in94_52 sn94_52 202000.000000
Rwneg94_53 in94_53 sn94_53 78000.000000
Rwneg94_54 in94_54 sn94_54 78000.000000
Rwneg94_55 in94_55 sn94_55 202000.000000
Rwneg94_56 in94_56 sn94_56 202000.000000
Rwneg94_57 in94_57 sn94_57 202000.000000
Rwneg94_58 in94_58 sn94_58 78000.000000
Rwneg94_59 in94_59 sn94_59 202000.000000
Rwneg94_60 in94_60 sn94_60 202000.000000
Rwneg94_61 in94_61 sn94_61 202000.000000
Rwneg94_62 in94_62 sn94_62 78000.000000
Rwneg94_63 in94_63 sn94_63 202000.000000
Rwneg94_64 in94_64 sn94_64 202000.000000
Rwneg94_65 in94_65 sn94_65 202000.000000
Rwneg94_66 in94_66 sn94_66 78000.000000
Rwneg94_67 in94_67 sn94_67 202000.000000
Rwneg94_68 in94_68 sn94_68 202000.000000
Rwneg94_69 in94_69 sn94_69 202000.000000
Rwneg94_70 in94_70 sn94_70 202000.000000
Rwneg94_71 in94_71 sn94_71 202000.000000
Rwneg94_72 in94_72 sn94_72 78000.000000
Rwneg94_73 in94_73 sn94_73 202000.000000
Rwneg94_74 in94_74 sn94_74 202000.000000
Rwneg94_75 in94_75 sn94_75 202000.000000
Rwneg94_76 in94_76 sn94_76 202000.000000
Rwneg94_77 in94_77 sn94_77 202000.000000
Rwneg94_78 in94_78 sn94_78 202000.000000
Rwneg94_79 in94_79 sn94_79 202000.000000
Rwneg94_80 in94_80 sn94_80 78000.000000
Rwneg94_81 in94_81 sn94_81 78000.000000
Rwneg94_82 in94_82 sn94_82 202000.000000
Rwneg94_83 in94_83 sn94_83 78000.000000
Rwneg94_84 in94_84 sn94_84 78000.000000
Rwneg95_1 in95_1 sn95_1 78000.000000
Rwneg95_2 in95_2 sn95_2 202000.000000
Rwneg95_3 in95_3 sn95_3 202000.000000
Rwneg95_4 in95_4 sn95_4 202000.000000
Rwneg95_5 in95_5 sn95_5 78000.000000
Rwneg95_6 in95_6 sn95_6 78000.000000
Rwneg95_7 in95_7 sn95_7 202000.000000
Rwneg95_8 in95_8 sn95_8 202000.000000
Rwneg95_9 in95_9 sn95_9 202000.000000
Rwneg95_10 in95_10 sn95_10 78000.000000
Rwneg95_11 in95_11 sn95_11 78000.000000
Rwneg95_12 in95_12 sn95_12 202000.000000
Rwneg95_13 in95_13 sn95_13 202000.000000
Rwneg95_14 in95_14 sn95_14 78000.000000
Rwneg95_15 in95_15 sn95_15 202000.000000
Rwneg95_16 in95_16 sn95_16 202000.000000
Rwneg95_17 in95_17 sn95_17 78000.000000
Rwneg95_18 in95_18 sn95_18 202000.000000
Rwneg95_19 in95_19 sn95_19 78000.000000
Rwneg95_20 in95_20 sn95_20 202000.000000
Rwneg95_21 in95_21 sn95_21 202000.000000
Rwneg95_22 in95_22 sn95_22 202000.000000
Rwneg95_23 in95_23 sn95_23 78000.000000
Rwneg95_24 in95_24 sn95_24 202000.000000
Rwneg95_25 in95_25 sn95_25 78000.000000
Rwneg95_26 in95_26 sn95_26 202000.000000
Rwneg95_27 in95_27 sn95_27 202000.000000
Rwneg95_28 in95_28 sn95_28 202000.000000
Rwneg95_29 in95_29 sn95_29 202000.000000
Rwneg95_30 in95_30 sn95_30 78000.000000
Rwneg95_31 in95_31 sn95_31 78000.000000
Rwneg95_32 in95_32 sn95_32 78000.000000
Rwneg95_33 in95_33 sn95_33 202000.000000
Rwneg95_34 in95_34 sn95_34 202000.000000
Rwneg95_35 in95_35 sn95_35 202000.000000
Rwneg95_36 in95_36 sn95_36 78000.000000
Rwneg95_37 in95_37 sn95_37 202000.000000
Rwneg95_38 in95_38 sn95_38 202000.000000
Rwneg95_39 in95_39 sn95_39 78000.000000
Rwneg95_40 in95_40 sn95_40 78000.000000
Rwneg95_41 in95_41 sn95_41 78000.000000
Rwneg95_42 in95_42 sn95_42 202000.000000
Rwneg95_43 in95_43 sn95_43 78000.000000
Rwneg95_44 in95_44 sn95_44 78000.000000
Rwneg95_45 in95_45 sn95_45 78000.000000
Rwneg95_46 in95_46 sn95_46 202000.000000
Rwneg95_47 in95_47 sn95_47 78000.000000
Rwneg95_48 in95_48 sn95_48 78000.000000
Rwneg95_49 in95_49 sn95_49 202000.000000
Rwneg95_50 in95_50 sn95_50 202000.000000
Rwneg95_51 in95_51 sn95_51 202000.000000
Rwneg95_52 in95_52 sn95_52 202000.000000
Rwneg95_53 in95_53 sn95_53 202000.000000
Rwneg95_54 in95_54 sn95_54 78000.000000
Rwneg95_55 in95_55 sn95_55 78000.000000
Rwneg95_56 in95_56 sn95_56 202000.000000
Rwneg95_57 in95_57 sn95_57 202000.000000
Rwneg95_58 in95_58 sn95_58 78000.000000
Rwneg95_59 in95_59 sn95_59 202000.000000
Rwneg95_60 in95_60 sn95_60 202000.000000
Rwneg95_61 in95_61 sn95_61 202000.000000
Rwneg95_62 in95_62 sn95_62 78000.000000
Rwneg95_63 in95_63 sn95_63 202000.000000
Rwneg95_64 in95_64 sn95_64 202000.000000
Rwneg95_65 in95_65 sn95_65 202000.000000
Rwneg95_66 in95_66 sn95_66 202000.000000
Rwneg95_67 in95_67 sn95_67 78000.000000
Rwneg95_68 in95_68 sn95_68 78000.000000
Rwneg95_69 in95_69 sn95_69 202000.000000
Rwneg95_70 in95_70 sn95_70 202000.000000
Rwneg95_71 in95_71 sn95_71 202000.000000
Rwneg95_72 in95_72 sn95_72 202000.000000
Rwneg95_73 in95_73 sn95_73 78000.000000
Rwneg95_74 in95_74 sn95_74 202000.000000
Rwneg95_75 in95_75 sn95_75 202000.000000
Rwneg95_76 in95_76 sn95_76 78000.000000
Rwneg95_77 in95_77 sn95_77 78000.000000
Rwneg95_78 in95_78 sn95_78 202000.000000
Rwneg95_79 in95_79 sn95_79 78000.000000
Rwneg95_80 in95_80 sn95_80 202000.000000
Rwneg95_81 in95_81 sn95_81 78000.000000
Rwneg95_82 in95_82 sn95_82 202000.000000
Rwneg95_83 in95_83 sn95_83 78000.000000
Rwneg95_84 in95_84 sn95_84 78000.000000
Rwneg96_1 in96_1 sn96_1 202000.000000
Rwneg96_2 in96_2 sn96_2 202000.000000
Rwneg96_3 in96_3 sn96_3 202000.000000
Rwneg96_4 in96_4 sn96_4 78000.000000
Rwneg96_5 in96_5 sn96_5 202000.000000
Rwneg96_6 in96_6 sn96_6 202000.000000
Rwneg96_7 in96_7 sn96_7 202000.000000
Rwneg96_8 in96_8 sn96_8 78000.000000
Rwneg96_9 in96_9 sn96_9 78000.000000
Rwneg96_10 in96_10 sn96_10 78000.000000
Rwneg96_11 in96_11 sn96_11 78000.000000
Rwneg96_12 in96_12 sn96_12 78000.000000
Rwneg96_13 in96_13 sn96_13 202000.000000
Rwneg96_14 in96_14 sn96_14 202000.000000
Rwneg96_15 in96_15 sn96_15 202000.000000
Rwneg96_16 in96_16 sn96_16 78000.000000
Rwneg96_17 in96_17 sn96_17 78000.000000
Rwneg96_18 in96_18 sn96_18 78000.000000
Rwneg96_19 in96_19 sn96_19 202000.000000
Rwneg96_20 in96_20 sn96_20 78000.000000
Rwneg96_21 in96_21 sn96_21 202000.000000
Rwneg96_22 in96_22 sn96_22 202000.000000
Rwneg96_23 in96_23 sn96_23 78000.000000
Rwneg96_24 in96_24 sn96_24 202000.000000
Rwneg96_25 in96_25 sn96_25 78000.000000
Rwneg96_26 in96_26 sn96_26 202000.000000
Rwneg96_27 in96_27 sn96_27 202000.000000
Rwneg96_28 in96_28 sn96_28 202000.000000
Rwneg96_29 in96_29 sn96_29 202000.000000
Rwneg96_30 in96_30 sn96_30 78000.000000
Rwneg96_31 in96_31 sn96_31 78000.000000
Rwneg96_32 in96_32 sn96_32 78000.000000
Rwneg96_33 in96_33 sn96_33 202000.000000
Rwneg96_34 in96_34 sn96_34 78000.000000
Rwneg96_35 in96_35 sn96_35 202000.000000
Rwneg96_36 in96_36 sn96_36 78000.000000
Rwneg96_37 in96_37 sn96_37 78000.000000
Rwneg96_38 in96_38 sn96_38 202000.000000
Rwneg96_39 in96_39 sn96_39 202000.000000
Rwneg96_40 in96_40 sn96_40 202000.000000
Rwneg96_41 in96_41 sn96_41 202000.000000
Rwneg96_42 in96_42 sn96_42 202000.000000
Rwneg96_43 in96_43 sn96_43 78000.000000
Rwneg96_44 in96_44 sn96_44 202000.000000
Rwneg96_45 in96_45 sn96_45 78000.000000
Rwneg96_46 in96_46 sn96_46 78000.000000
Rwneg96_47 in96_47 sn96_47 202000.000000
Rwneg96_48 in96_48 sn96_48 202000.000000
Rwneg96_49 in96_49 sn96_49 202000.000000
Rwneg96_50 in96_50 sn96_50 202000.000000
Rwneg96_51 in96_51 sn96_51 202000.000000
Rwneg96_52 in96_52 sn96_52 202000.000000
Rwneg96_53 in96_53 sn96_53 78000.000000
Rwneg96_54 in96_54 sn96_54 202000.000000
Rwneg96_55 in96_55 sn96_55 202000.000000
Rwneg96_56 in96_56 sn96_56 78000.000000
Rwneg96_57 in96_57 sn96_57 202000.000000
Rwneg96_58 in96_58 sn96_58 78000.000000
Rwneg96_59 in96_59 sn96_59 78000.000000
Rwneg96_60 in96_60 sn96_60 202000.000000
Rwneg96_61 in96_61 sn96_61 78000.000000
Rwneg96_62 in96_62 sn96_62 78000.000000
Rwneg96_63 in96_63 sn96_63 78000.000000
Rwneg96_64 in96_64 sn96_64 202000.000000
Rwneg96_65 in96_65 sn96_65 202000.000000
Rwneg96_66 in96_66 sn96_66 78000.000000
Rwneg96_67 in96_67 sn96_67 202000.000000
Rwneg96_68 in96_68 sn96_68 78000.000000
Rwneg96_69 in96_69 sn96_69 78000.000000
Rwneg96_70 in96_70 sn96_70 78000.000000
Rwneg96_71 in96_71 sn96_71 78000.000000
Rwneg96_72 in96_72 sn96_72 202000.000000
Rwneg96_73 in96_73 sn96_73 78000.000000
Rwneg96_74 in96_74 sn96_74 202000.000000
Rwneg96_75 in96_75 sn96_75 202000.000000
Rwneg96_76 in96_76 sn96_76 202000.000000
Rwneg96_77 in96_77 sn96_77 78000.000000
Rwneg96_78 in96_78 sn96_78 202000.000000
Rwneg96_79 in96_79 sn96_79 78000.000000
Rwneg96_80 in96_80 sn96_80 78000.000000
Rwneg96_81 in96_81 sn96_81 202000.000000
Rwneg96_82 in96_82 sn96_82 78000.000000
Rwneg96_83 in96_83 sn96_83 202000.000000
Rwneg96_84 in96_84 sn96_84 202000.000000
Rwneg97_1 in97_1 sn97_1 78000.000000
Rwneg97_2 in97_2 sn97_2 202000.000000
Rwneg97_3 in97_3 sn97_3 78000.000000
Rwneg97_4 in97_4 sn97_4 202000.000000
Rwneg97_5 in97_5 sn97_5 78000.000000
Rwneg97_6 in97_6 sn97_6 202000.000000
Rwneg97_7 in97_7 sn97_7 202000.000000
Rwneg97_8 in97_8 sn97_8 202000.000000
Rwneg97_9 in97_9 sn97_9 202000.000000
Rwneg97_10 in97_10 sn97_10 78000.000000
Rwneg97_11 in97_11 sn97_11 78000.000000
Rwneg97_12 in97_12 sn97_12 202000.000000
Rwneg97_13 in97_13 sn97_13 78000.000000
Rwneg97_14 in97_14 sn97_14 78000.000000
Rwneg97_15 in97_15 sn97_15 202000.000000
Rwneg97_16 in97_16 sn97_16 202000.000000
Rwneg97_17 in97_17 sn97_17 202000.000000
Rwneg97_18 in97_18 sn97_18 78000.000000
Rwneg97_19 in97_19 sn97_19 202000.000000
Rwneg97_20 in97_20 sn97_20 78000.000000
Rwneg97_21 in97_21 sn97_21 202000.000000
Rwneg97_22 in97_22 sn97_22 202000.000000
Rwneg97_23 in97_23 sn97_23 202000.000000
Rwneg97_24 in97_24 sn97_24 78000.000000
Rwneg97_25 in97_25 sn97_25 202000.000000
Rwneg97_26 in97_26 sn97_26 202000.000000
Rwneg97_27 in97_27 sn97_27 202000.000000
Rwneg97_28 in97_28 sn97_28 78000.000000
Rwneg97_29 in97_29 sn97_29 78000.000000
Rwneg97_30 in97_30 sn97_30 202000.000000
Rwneg97_31 in97_31 sn97_31 202000.000000
Rwneg97_32 in97_32 sn97_32 78000.000000
Rwneg97_33 in97_33 sn97_33 78000.000000
Rwneg97_34 in97_34 sn97_34 78000.000000
Rwneg97_35 in97_35 sn97_35 78000.000000
Rwneg97_36 in97_36 sn97_36 78000.000000
Rwneg97_37 in97_37 sn97_37 78000.000000
Rwneg97_38 in97_38 sn97_38 78000.000000
Rwneg97_39 in97_39 sn97_39 78000.000000
Rwneg97_40 in97_40 sn97_40 78000.000000
Rwneg97_41 in97_41 sn97_41 202000.000000
Rwneg97_42 in97_42 sn97_42 78000.000000
Rwneg97_43 in97_43 sn97_43 202000.000000
Rwneg97_44 in97_44 sn97_44 202000.000000
Rwneg97_45 in97_45 sn97_45 202000.000000
Rwneg97_46 in97_46 sn97_46 78000.000000
Rwneg97_47 in97_47 sn97_47 78000.000000
Rwneg97_48 in97_48 sn97_48 78000.000000
Rwneg97_49 in97_49 sn97_49 202000.000000
Rwneg97_50 in97_50 sn97_50 78000.000000
Rwneg97_51 in97_51 sn97_51 78000.000000
Rwneg97_52 in97_52 sn97_52 202000.000000
Rwneg97_53 in97_53 sn97_53 78000.000000
Rwneg97_54 in97_54 sn97_54 202000.000000
Rwneg97_55 in97_55 sn97_55 78000.000000
Rwneg97_56 in97_56 sn97_56 202000.000000
Rwneg97_57 in97_57 sn97_57 78000.000000
Rwneg97_58 in97_58 sn97_58 202000.000000
Rwneg97_59 in97_59 sn97_59 78000.000000
Rwneg97_60 in97_60 sn97_60 202000.000000
Rwneg97_61 in97_61 sn97_61 202000.000000
Rwneg97_62 in97_62 sn97_62 78000.000000
Rwneg97_63 in97_63 sn97_63 202000.000000
Rwneg97_64 in97_64 sn97_64 78000.000000
Rwneg97_65 in97_65 sn97_65 202000.000000
Rwneg97_66 in97_66 sn97_66 202000.000000
Rwneg97_67 in97_67 sn97_67 78000.000000
Rwneg97_68 in97_68 sn97_68 202000.000000
Rwneg97_69 in97_69 sn97_69 202000.000000
Rwneg97_70 in97_70 sn97_70 202000.000000
Rwneg97_71 in97_71 sn97_71 202000.000000
Rwneg97_72 in97_72 sn97_72 202000.000000
Rwneg97_73 in97_73 sn97_73 202000.000000
Rwneg97_74 in97_74 sn97_74 202000.000000
Rwneg97_75 in97_75 sn97_75 78000.000000
Rwneg97_76 in97_76 sn97_76 202000.000000
Rwneg97_77 in97_77 sn97_77 202000.000000
Rwneg97_78 in97_78 sn97_78 202000.000000
Rwneg97_79 in97_79 sn97_79 202000.000000
Rwneg97_80 in97_80 sn97_80 78000.000000
Rwneg97_81 in97_81 sn97_81 202000.000000
Rwneg97_82 in97_82 sn97_82 202000.000000
Rwneg97_83 in97_83 sn97_83 202000.000000
Rwneg97_84 in97_84 sn97_84 202000.000000
Rwneg98_1 in98_1 sn98_1 202000.000000
Rwneg98_2 in98_2 sn98_2 202000.000000
Rwneg98_3 in98_3 sn98_3 202000.000000
Rwneg98_4 in98_4 sn98_4 202000.000000
Rwneg98_5 in98_5 sn98_5 202000.000000
Rwneg98_6 in98_6 sn98_6 78000.000000
Rwneg98_7 in98_7 sn98_7 78000.000000
Rwneg98_8 in98_8 sn98_8 202000.000000
Rwneg98_9 in98_9 sn98_9 202000.000000
Rwneg98_10 in98_10 sn98_10 202000.000000
Rwneg98_11 in98_11 sn98_11 202000.000000
Rwneg98_12 in98_12 sn98_12 202000.000000
Rwneg98_13 in98_13 sn98_13 202000.000000
Rwneg98_14 in98_14 sn98_14 78000.000000
Rwneg98_15 in98_15 sn98_15 78000.000000
Rwneg98_16 in98_16 sn98_16 78000.000000
Rwneg98_17 in98_17 sn98_17 202000.000000
Rwneg98_18 in98_18 sn98_18 202000.000000
Rwneg98_19 in98_19 sn98_19 78000.000000
Rwneg98_20 in98_20 sn98_20 78000.000000
Rwneg98_21 in98_21 sn98_21 78000.000000
Rwneg98_22 in98_22 sn98_22 78000.000000
Rwneg98_23 in98_23 sn98_23 78000.000000
Rwneg98_24 in98_24 sn98_24 202000.000000
Rwneg98_25 in98_25 sn98_25 202000.000000
Rwneg98_26 in98_26 sn98_26 202000.000000
Rwneg98_27 in98_27 sn98_27 202000.000000
Rwneg98_28 in98_28 sn98_28 78000.000000
Rwneg98_29 in98_29 sn98_29 78000.000000
Rwneg98_30 in98_30 sn98_30 202000.000000
Rwneg98_31 in98_31 sn98_31 78000.000000
Rwneg98_32 in98_32 sn98_32 202000.000000
Rwneg98_33 in98_33 sn98_33 78000.000000
Rwneg98_34 in98_34 sn98_34 202000.000000
Rwneg98_35 in98_35 sn98_35 78000.000000
Rwneg98_36 in98_36 sn98_36 202000.000000
Rwneg98_37 in98_37 sn98_37 78000.000000
Rwneg98_38 in98_38 sn98_38 78000.000000
Rwneg98_39 in98_39 sn98_39 78000.000000
Rwneg98_40 in98_40 sn98_40 78000.000000
Rwneg98_41 in98_41 sn98_41 78000.000000
Rwneg98_42 in98_42 sn98_42 78000.000000
Rwneg98_43 in98_43 sn98_43 78000.000000
Rwneg98_44 in98_44 sn98_44 202000.000000
Rwneg98_45 in98_45 sn98_45 78000.000000
Rwneg98_46 in98_46 sn98_46 78000.000000
Rwneg98_47 in98_47 sn98_47 202000.000000
Rwneg98_48 in98_48 sn98_48 202000.000000
Rwneg98_49 in98_49 sn98_49 202000.000000
Rwneg98_50 in98_50 sn98_50 78000.000000
Rwneg98_51 in98_51 sn98_51 78000.000000
Rwneg98_52 in98_52 sn98_52 78000.000000
Rwneg98_53 in98_53 sn98_53 78000.000000
Rwneg98_54 in98_54 sn98_54 78000.000000
Rwneg98_55 in98_55 sn98_55 78000.000000
Rwneg98_56 in98_56 sn98_56 202000.000000
Rwneg98_57 in98_57 sn98_57 202000.000000
Rwneg98_58 in98_58 sn98_58 78000.000000
Rwneg98_59 in98_59 sn98_59 202000.000000
Rwneg98_60 in98_60 sn98_60 202000.000000
Rwneg98_61 in98_61 sn98_61 78000.000000
Rwneg98_62 in98_62 sn98_62 202000.000000
Rwneg98_63 in98_63 sn98_63 202000.000000
Rwneg98_64 in98_64 sn98_64 202000.000000
Rwneg98_65 in98_65 sn98_65 78000.000000
Rwneg98_66 in98_66 sn98_66 202000.000000
Rwneg98_67 in98_67 sn98_67 78000.000000
Rwneg98_68 in98_68 sn98_68 202000.000000
Rwneg98_69 in98_69 sn98_69 202000.000000
Rwneg98_70 in98_70 sn98_70 202000.000000
Rwneg98_71 in98_71 sn98_71 202000.000000
Rwneg98_72 in98_72 sn98_72 202000.000000
Rwneg98_73 in98_73 sn98_73 202000.000000
Rwneg98_74 in98_74 sn98_74 202000.000000
Rwneg98_75 in98_75 sn98_75 78000.000000
Rwneg98_76 in98_76 sn98_76 202000.000000
Rwneg98_77 in98_77 sn98_77 78000.000000
Rwneg98_78 in98_78 sn98_78 202000.000000
Rwneg98_79 in98_79 sn98_79 202000.000000
Rwneg98_80 in98_80 sn98_80 78000.000000
Rwneg98_81 in98_81 sn98_81 202000.000000
Rwneg98_82 in98_82 sn98_82 202000.000000
Rwneg98_83 in98_83 sn98_83 78000.000000
Rwneg98_84 in98_84 sn98_84 78000.000000
Rwneg99_1 in99_1 sn99_1 202000.000000
Rwneg99_2 in99_2 sn99_2 202000.000000
Rwneg99_3 in99_3 sn99_3 78000.000000
Rwneg99_4 in99_4 sn99_4 202000.000000
Rwneg99_5 in99_5 sn99_5 202000.000000
Rwneg99_6 in99_6 sn99_6 202000.000000
Rwneg99_7 in99_7 sn99_7 78000.000000
Rwneg99_8 in99_8 sn99_8 78000.000000
Rwneg99_9 in99_9 sn99_9 202000.000000
Rwneg99_10 in99_10 sn99_10 202000.000000
Rwneg99_11 in99_11 sn99_11 202000.000000
Rwneg99_12 in99_12 sn99_12 202000.000000
Rwneg99_13 in99_13 sn99_13 202000.000000
Rwneg99_14 in99_14 sn99_14 202000.000000
Rwneg99_15 in99_15 sn99_15 78000.000000
Rwneg99_16 in99_16 sn99_16 202000.000000
Rwneg99_17 in99_17 sn99_17 202000.000000
Rwneg99_18 in99_18 sn99_18 202000.000000
Rwneg99_19 in99_19 sn99_19 202000.000000
Rwneg99_20 in99_20 sn99_20 78000.000000
Rwneg99_21 in99_21 sn99_21 202000.000000
Rwneg99_22 in99_22 sn99_22 202000.000000
Rwneg99_23 in99_23 sn99_23 202000.000000
Rwneg99_24 in99_24 sn99_24 78000.000000
Rwneg99_25 in99_25 sn99_25 202000.000000
Rwneg99_26 in99_26 sn99_26 202000.000000
Rwneg99_27 in99_27 sn99_27 202000.000000
Rwneg99_28 in99_28 sn99_28 202000.000000
Rwneg99_29 in99_29 sn99_29 202000.000000
Rwneg99_30 in99_30 sn99_30 78000.000000
Rwneg99_31 in99_31 sn99_31 202000.000000
Rwneg99_32 in99_32 sn99_32 202000.000000
Rwneg99_33 in99_33 sn99_33 78000.000000
Rwneg99_34 in99_34 sn99_34 202000.000000
Rwneg99_35 in99_35 sn99_35 78000.000000
Rwneg99_36 in99_36 sn99_36 78000.000000
Rwneg99_37 in99_37 sn99_37 78000.000000
Rwneg99_38 in99_38 sn99_38 78000.000000
Rwneg99_39 in99_39 sn99_39 202000.000000
Rwneg99_40 in99_40 sn99_40 202000.000000
Rwneg99_41 in99_41 sn99_41 78000.000000
Rwneg99_42 in99_42 sn99_42 78000.000000
Rwneg99_43 in99_43 sn99_43 78000.000000
Rwneg99_44 in99_44 sn99_44 202000.000000
Rwneg99_45 in99_45 sn99_45 202000.000000
Rwneg99_46 in99_46 sn99_46 202000.000000
Rwneg99_47 in99_47 sn99_47 202000.000000
Rwneg99_48 in99_48 sn99_48 78000.000000
Rwneg99_49 in99_49 sn99_49 78000.000000
Rwneg99_50 in99_50 sn99_50 78000.000000
Rwneg99_51 in99_51 sn99_51 202000.000000
Rwneg99_52 in99_52 sn99_52 78000.000000
Rwneg99_53 in99_53 sn99_53 202000.000000
Rwneg99_54 in99_54 sn99_54 202000.000000
Rwneg99_55 in99_55 sn99_55 78000.000000
Rwneg99_56 in99_56 sn99_56 202000.000000
Rwneg99_57 in99_57 sn99_57 78000.000000
Rwneg99_58 in99_58 sn99_58 202000.000000
Rwneg99_59 in99_59 sn99_59 78000.000000
Rwneg99_60 in99_60 sn99_60 202000.000000
Rwneg99_61 in99_61 sn99_61 202000.000000
Rwneg99_62 in99_62 sn99_62 202000.000000
Rwneg99_63 in99_63 sn99_63 78000.000000
Rwneg99_64 in99_64 sn99_64 78000.000000
Rwneg99_65 in99_65 sn99_65 78000.000000
Rwneg99_66 in99_66 sn99_66 78000.000000
Rwneg99_67 in99_67 sn99_67 202000.000000
Rwneg99_68 in99_68 sn99_68 202000.000000
Rwneg99_69 in99_69 sn99_69 202000.000000
Rwneg99_70 in99_70 sn99_70 78000.000000
Rwneg99_71 in99_71 sn99_71 202000.000000
Rwneg99_72 in99_72 sn99_72 78000.000000
Rwneg99_73 in99_73 sn99_73 202000.000000
Rwneg99_74 in99_74 sn99_74 202000.000000
Rwneg99_75 in99_75 sn99_75 78000.000000
Rwneg99_76 in99_76 sn99_76 78000.000000
Rwneg99_77 in99_77 sn99_77 202000.000000
Rwneg99_78 in99_78 sn99_78 202000.000000
Rwneg99_79 in99_79 sn99_79 202000.000000
Rwneg99_80 in99_80 sn99_80 202000.000000
Rwneg99_81 in99_81 sn99_81 202000.000000
Rwneg99_82 in99_82 sn99_82 202000.000000
Rwneg99_83 in99_83 sn99_83 202000.000000
Rwneg99_84 in99_84 sn99_84 78000.000000
Rwneg100_1 in100_1 sn100_1 202000.000000
Rwneg100_2 in100_2 sn100_2 202000.000000
Rwneg100_3 in100_3 sn100_3 78000.000000
Rwneg100_4 in100_4 sn100_4 78000.000000
Rwneg100_5 in100_5 sn100_5 78000.000000
Rwneg100_6 in100_6 sn100_6 202000.000000
Rwneg100_7 in100_7 sn100_7 78000.000000
Rwneg100_8 in100_8 sn100_8 78000.000000
Rwneg100_9 in100_9 sn100_9 78000.000000
Rwneg100_10 in100_10 sn100_10 78000.000000
Rwneg100_11 in100_11 sn100_11 202000.000000
Rwneg100_12 in100_12 sn100_12 202000.000000
Rwneg100_13 in100_13 sn100_13 78000.000000
Rwneg100_14 in100_14 sn100_14 78000.000000
Rwneg100_15 in100_15 sn100_15 202000.000000
Rwneg100_16 in100_16 sn100_16 202000.000000
Rwneg100_17 in100_17 sn100_17 202000.000000
Rwneg100_18 in100_18 sn100_18 202000.000000
Rwneg100_19 in100_19 sn100_19 202000.000000
Rwneg100_20 in100_20 sn100_20 202000.000000
Rwneg100_21 in100_21 sn100_21 202000.000000
Rwneg100_22 in100_22 sn100_22 78000.000000
Rwneg100_23 in100_23 sn100_23 202000.000000
Rwneg100_24 in100_24 sn100_24 78000.000000
Rwneg100_25 in100_25 sn100_25 78000.000000
Rwneg100_26 in100_26 sn100_26 78000.000000
Rwneg100_27 in100_27 sn100_27 78000.000000
Rwneg100_28 in100_28 sn100_28 202000.000000
Rwneg100_29 in100_29 sn100_29 78000.000000
Rwneg100_30 in100_30 sn100_30 202000.000000
Rwneg100_31 in100_31 sn100_31 78000.000000
Rwneg100_32 in100_32 sn100_32 202000.000000
Rwneg100_33 in100_33 sn100_33 202000.000000
Rwneg100_34 in100_34 sn100_34 78000.000000
Rwneg100_35 in100_35 sn100_35 78000.000000
Rwneg100_36 in100_36 sn100_36 78000.000000
Rwneg100_37 in100_37 sn100_37 202000.000000
Rwneg100_38 in100_38 sn100_38 202000.000000
Rwneg100_39 in100_39 sn100_39 78000.000000
Rwneg100_40 in100_40 sn100_40 202000.000000
Rwneg100_41 in100_41 sn100_41 78000.000000
Rwneg100_42 in100_42 sn100_42 202000.000000
Rwneg100_43 in100_43 sn100_43 202000.000000
Rwneg100_44 in100_44 sn100_44 78000.000000
Rwneg100_45 in100_45 sn100_45 202000.000000
Rwneg100_46 in100_46 sn100_46 202000.000000
Rwneg100_47 in100_47 sn100_47 78000.000000
Rwneg100_48 in100_48 sn100_48 78000.000000
Rwneg100_49 in100_49 sn100_49 202000.000000
Rwneg100_50 in100_50 sn100_50 78000.000000
Rwneg100_51 in100_51 sn100_51 78000.000000
Rwneg100_52 in100_52 sn100_52 202000.000000
Rwneg100_53 in100_53 sn100_53 202000.000000
Rwneg100_54 in100_54 sn100_54 202000.000000
Rwneg100_55 in100_55 sn100_55 202000.000000
Rwneg100_56 in100_56 sn100_56 202000.000000
Rwneg100_57 in100_57 sn100_57 78000.000000
Rwneg100_58 in100_58 sn100_58 202000.000000
Rwneg100_59 in100_59 sn100_59 202000.000000
Rwneg100_60 in100_60 sn100_60 78000.000000
Rwneg100_61 in100_61 sn100_61 202000.000000
Rwneg100_62 in100_62 sn100_62 78000.000000
Rwneg100_63 in100_63 sn100_63 202000.000000
Rwneg100_64 in100_64 sn100_64 202000.000000
Rwneg100_65 in100_65 sn100_65 78000.000000
Rwneg100_66 in100_66 sn100_66 78000.000000
Rwneg100_67 in100_67 sn100_67 78000.000000
Rwneg100_68 in100_68 sn100_68 202000.000000
Rwneg100_69 in100_69 sn100_69 202000.000000
Rwneg100_70 in100_70 sn100_70 78000.000000
Rwneg100_71 in100_71 sn100_71 202000.000000
Rwneg100_72 in100_72 sn100_72 78000.000000
Rwneg100_73 in100_73 sn100_73 202000.000000
Rwneg100_74 in100_74 sn100_74 78000.000000
Rwneg100_75 in100_75 sn100_75 78000.000000
Rwneg100_76 in100_76 sn100_76 78000.000000
Rwneg100_77 in100_77 sn100_77 202000.000000
Rwneg100_78 in100_78 sn100_78 78000.000000
Rwneg100_79 in100_79 sn100_79 202000.000000
Rwneg100_80 in100_80 sn100_80 202000.000000
Rwneg100_81 in100_81 sn100_81 202000.000000
Rwneg100_82 in100_82 sn100_82 78000.000000
Rwneg100_83 in100_83 sn100_83 202000.000000
Rwneg100_84 in100_84 sn100_84 202000.000000
Rwneg101_1 in101_1 sn101_1 202000.000000
Rwneg101_2 in101_2 sn101_2 202000.000000
Rwneg101_3 in101_3 sn101_3 78000.000000
Rwneg101_4 in101_4 sn101_4 78000.000000
Rwneg101_5 in101_5 sn101_5 78000.000000
Rwneg101_6 in101_6 sn101_6 202000.000000
Rwneg101_7 in101_7 sn101_7 202000.000000
Rwneg101_8 in101_8 sn101_8 202000.000000
Rwneg101_9 in101_9 sn101_9 78000.000000
Rwneg101_10 in101_10 sn101_10 202000.000000
Rwneg101_11 in101_11 sn101_11 202000.000000
Rwneg101_12 in101_12 sn101_12 78000.000000
Rwneg101_13 in101_13 sn101_13 202000.000000
Rwneg101_14 in101_14 sn101_14 202000.000000
Rwneg101_15 in101_15 sn101_15 202000.000000
Rwneg101_16 in101_16 sn101_16 78000.000000
Rwneg101_17 in101_17 sn101_17 78000.000000
Rwneg101_18 in101_18 sn101_18 78000.000000
Rwneg101_19 in101_19 sn101_19 202000.000000
Rwneg101_20 in101_20 sn101_20 202000.000000
Rwneg101_21 in101_21 sn101_21 202000.000000
Rwneg101_22 in101_22 sn101_22 78000.000000
Rwneg101_23 in101_23 sn101_23 202000.000000
Rwneg101_24 in101_24 sn101_24 202000.000000
Rwneg101_25 in101_25 sn101_25 202000.000000
Rwneg101_26 in101_26 sn101_26 78000.000000
Rwneg101_27 in101_27 sn101_27 78000.000000
Rwneg101_28 in101_28 sn101_28 202000.000000
Rwneg101_29 in101_29 sn101_29 78000.000000
Rwneg101_30 in101_30 sn101_30 202000.000000
Rwneg101_31 in101_31 sn101_31 78000.000000
Rwneg101_32 in101_32 sn101_32 78000.000000
Rwneg101_33 in101_33 sn101_33 78000.000000
Rwneg101_34 in101_34 sn101_34 202000.000000
Rwneg101_35 in101_35 sn101_35 78000.000000
Rwneg101_36 in101_36 sn101_36 202000.000000
Rwneg101_37 in101_37 sn101_37 202000.000000
Rwneg101_38 in101_38 sn101_38 202000.000000
Rwneg101_39 in101_39 sn101_39 202000.000000
Rwneg101_40 in101_40 sn101_40 78000.000000
Rwneg101_41 in101_41 sn101_41 78000.000000
Rwneg101_42 in101_42 sn101_42 202000.000000
Rwneg101_43 in101_43 sn101_43 78000.000000
Rwneg101_44 in101_44 sn101_44 202000.000000
Rwneg101_45 in101_45 sn101_45 202000.000000
Rwneg101_46 in101_46 sn101_46 202000.000000
Rwneg101_47 in101_47 sn101_47 202000.000000
Rwneg101_48 in101_48 sn101_48 202000.000000
Rwneg101_49 in101_49 sn101_49 202000.000000
Rwneg101_50 in101_50 sn101_50 202000.000000
Rwneg101_51 in101_51 sn101_51 78000.000000
Rwneg101_52 in101_52 sn101_52 202000.000000
Rwneg101_53 in101_53 sn101_53 202000.000000
Rwneg101_54 in101_54 sn101_54 78000.000000
Rwneg101_55 in101_55 sn101_55 78000.000000
Rwneg101_56 in101_56 sn101_56 202000.000000
Rwneg101_57 in101_57 sn101_57 78000.000000
Rwneg101_58 in101_58 sn101_58 202000.000000
Rwneg101_59 in101_59 sn101_59 202000.000000
Rwneg101_60 in101_60 sn101_60 202000.000000
Rwneg101_61 in101_61 sn101_61 78000.000000
Rwneg101_62 in101_62 sn101_62 78000.000000
Rwneg101_63 in101_63 sn101_63 202000.000000
Rwneg101_64 in101_64 sn101_64 78000.000000
Rwneg101_65 in101_65 sn101_65 202000.000000
Rwneg101_66 in101_66 sn101_66 78000.000000
Rwneg101_67 in101_67 sn101_67 202000.000000
Rwneg101_68 in101_68 sn101_68 78000.000000
Rwneg101_69 in101_69 sn101_69 78000.000000
Rwneg101_70 in101_70 sn101_70 78000.000000
Rwneg101_71 in101_71 sn101_71 202000.000000
Rwneg101_72 in101_72 sn101_72 78000.000000
Rwneg101_73 in101_73 sn101_73 78000.000000
Rwneg101_74 in101_74 sn101_74 78000.000000
Rwneg101_75 in101_75 sn101_75 202000.000000
Rwneg101_76 in101_76 sn101_76 202000.000000
Rwneg101_77 in101_77 sn101_77 202000.000000
Rwneg101_78 in101_78 sn101_78 78000.000000
Rwneg101_79 in101_79 sn101_79 202000.000000
Rwneg101_80 in101_80 sn101_80 78000.000000
Rwneg101_81 in101_81 sn101_81 202000.000000
Rwneg101_82 in101_82 sn101_82 202000.000000
Rwneg101_83 in101_83 sn101_83 78000.000000
Rwneg101_84 in101_84 sn101_84 202000.000000
Rwneg102_1 in102_1 sn102_1 78000.000000
Rwneg102_2 in102_2 sn102_2 202000.000000
Rwneg102_3 in102_3 sn102_3 78000.000000
Rwneg102_4 in102_4 sn102_4 202000.000000
Rwneg102_5 in102_5 sn102_5 78000.000000
Rwneg102_6 in102_6 sn102_6 202000.000000
Rwneg102_7 in102_7 sn102_7 202000.000000
Rwneg102_8 in102_8 sn102_8 202000.000000
Rwneg102_9 in102_9 sn102_9 202000.000000
Rwneg102_10 in102_10 sn102_10 202000.000000
Rwneg102_11 in102_11 sn102_11 202000.000000
Rwneg102_12 in102_12 sn102_12 78000.000000
Rwneg102_13 in102_13 sn102_13 202000.000000
Rwneg102_14 in102_14 sn102_14 78000.000000
Rwneg102_15 in102_15 sn102_15 202000.000000
Rwneg102_16 in102_16 sn102_16 78000.000000
Rwneg102_17 in102_17 sn102_17 202000.000000
Rwneg102_18 in102_18 sn102_18 78000.000000
Rwneg102_19 in102_19 sn102_19 78000.000000
Rwneg102_20 in102_20 sn102_20 78000.000000
Rwneg102_21 in102_21 sn102_21 202000.000000
Rwneg102_22 in102_22 sn102_22 202000.000000
Rwneg102_23 in102_23 sn102_23 202000.000000
Rwneg102_24 in102_24 sn102_24 202000.000000
Rwneg102_25 in102_25 sn102_25 78000.000000
Rwneg102_26 in102_26 sn102_26 78000.000000
Rwneg102_27 in102_27 sn102_27 202000.000000
Rwneg102_28 in102_28 sn102_28 78000.000000
Rwneg102_29 in102_29 sn102_29 78000.000000
Rwneg102_30 in102_30 sn102_30 202000.000000
Rwneg102_31 in102_31 sn102_31 202000.000000
Rwneg102_32 in102_32 sn102_32 78000.000000
Rwneg102_33 in102_33 sn102_33 78000.000000
Rwneg102_34 in102_34 sn102_34 78000.000000
Rwneg102_35 in102_35 sn102_35 78000.000000
Rwneg102_36 in102_36 sn102_36 202000.000000
Rwneg102_37 in102_37 sn102_37 202000.000000
Rwneg102_38 in102_38 sn102_38 78000.000000
Rwneg102_39 in102_39 sn102_39 78000.000000
Rwneg102_40 in102_40 sn102_40 78000.000000
Rwneg102_41 in102_41 sn102_41 78000.000000
Rwneg102_42 in102_42 sn102_42 78000.000000
Rwneg102_43 in102_43 sn102_43 202000.000000
Rwneg102_44 in102_44 sn102_44 202000.000000
Rwneg102_45 in102_45 sn102_45 78000.000000
Rwneg102_46 in102_46 sn102_46 78000.000000
Rwneg102_47 in102_47 sn102_47 202000.000000
Rwneg102_48 in102_48 sn102_48 78000.000000
Rwneg102_49 in102_49 sn102_49 78000.000000
Rwneg102_50 in102_50 sn102_50 78000.000000
Rwneg102_51 in102_51 sn102_51 78000.000000
Rwneg102_52 in102_52 sn102_52 202000.000000
Rwneg102_53 in102_53 sn102_53 78000.000000
Rwneg102_54 in102_54 sn102_54 78000.000000
Rwneg102_55 in102_55 sn102_55 202000.000000
Rwneg102_56 in102_56 sn102_56 202000.000000
Rwneg102_57 in102_57 sn102_57 78000.000000
Rwneg102_58 in102_58 sn102_58 202000.000000
Rwneg102_59 in102_59 sn102_59 202000.000000
Rwneg102_60 in102_60 sn102_60 202000.000000
Rwneg102_61 in102_61 sn102_61 202000.000000
Rwneg102_62 in102_62 sn102_62 202000.000000
Rwneg102_63 in102_63 sn102_63 202000.000000
Rwneg102_64 in102_64 sn102_64 202000.000000
Rwneg102_65 in102_65 sn102_65 202000.000000
Rwneg102_66 in102_66 sn102_66 202000.000000
Rwneg102_67 in102_67 sn102_67 78000.000000
Rwneg102_68 in102_68 sn102_68 202000.000000
Rwneg102_69 in102_69 sn102_69 202000.000000
Rwneg102_70 in102_70 sn102_70 202000.000000
Rwneg102_71 in102_71 sn102_71 202000.000000
Rwneg102_72 in102_72 sn102_72 202000.000000
Rwneg102_73 in102_73 sn102_73 202000.000000
Rwneg102_74 in102_74 sn102_74 202000.000000
Rwneg102_75 in102_75 sn102_75 78000.000000
Rwneg102_76 in102_76 sn102_76 202000.000000
Rwneg102_77 in102_77 sn102_77 202000.000000
Rwneg102_78 in102_78 sn102_78 202000.000000
Rwneg102_79 in102_79 sn102_79 202000.000000
Rwneg102_80 in102_80 sn102_80 78000.000000
Rwneg102_81 in102_81 sn102_81 202000.000000
Rwneg102_82 in102_82 sn102_82 202000.000000
Rwneg102_83 in102_83 sn102_83 78000.000000
Rwneg102_84 in102_84 sn102_84 78000.000000
Rwneg103_1 in103_1 sn103_1 78000.000000
Rwneg103_2 in103_2 sn103_2 78000.000000
Rwneg103_3 in103_3 sn103_3 202000.000000
Rwneg103_4 in103_4 sn103_4 78000.000000
Rwneg103_5 in103_5 sn103_5 78000.000000
Rwneg103_6 in103_6 sn103_6 78000.000000
Rwneg103_7 in103_7 sn103_7 202000.000000
Rwneg103_8 in103_8 sn103_8 202000.000000
Rwneg103_9 in103_9 sn103_9 78000.000000
Rwneg103_10 in103_10 sn103_10 202000.000000
Rwneg103_11 in103_11 sn103_11 202000.000000
Rwneg103_12 in103_12 sn103_12 78000.000000
Rwneg103_13 in103_13 sn103_13 78000.000000
Rwneg103_14 in103_14 sn103_14 202000.000000
Rwneg103_15 in103_15 sn103_15 202000.000000
Rwneg103_16 in103_16 sn103_16 78000.000000
Rwneg103_17 in103_17 sn103_17 78000.000000
Rwneg103_18 in103_18 sn103_18 78000.000000
Rwneg103_19 in103_19 sn103_19 78000.000000
Rwneg103_20 in103_20 sn103_20 202000.000000
Rwneg103_21 in103_21 sn103_21 202000.000000
Rwneg103_22 in103_22 sn103_22 78000.000000
Rwneg103_23 in103_23 sn103_23 202000.000000
Rwneg103_24 in103_24 sn103_24 78000.000000
Rwneg103_25 in103_25 sn103_25 78000.000000
Rwneg103_26 in103_26 sn103_26 202000.000000
Rwneg103_27 in103_27 sn103_27 78000.000000
Rwneg103_28 in103_28 sn103_28 202000.000000
Rwneg103_29 in103_29 sn103_29 202000.000000
Rwneg103_30 in103_30 sn103_30 202000.000000
Rwneg103_31 in103_31 sn103_31 78000.000000
Rwneg103_32 in103_32 sn103_32 202000.000000
Rwneg103_33 in103_33 sn103_33 202000.000000
Rwneg103_34 in103_34 sn103_34 202000.000000
Rwneg103_35 in103_35 sn103_35 202000.000000
Rwneg103_36 in103_36 sn103_36 78000.000000
Rwneg103_37 in103_37 sn103_37 202000.000000
Rwneg103_38 in103_38 sn103_38 202000.000000
Rwneg103_39 in103_39 sn103_39 78000.000000
Rwneg103_40 in103_40 sn103_40 202000.000000
Rwneg103_41 in103_41 sn103_41 202000.000000
Rwneg103_42 in103_42 sn103_42 202000.000000
Rwneg103_43 in103_43 sn103_43 202000.000000
Rwneg103_44 in103_44 sn103_44 78000.000000
Rwneg103_45 in103_45 sn103_45 78000.000000
Rwneg103_46 in103_46 sn103_46 202000.000000
Rwneg103_47 in103_47 sn103_47 78000.000000
Rwneg103_48 in103_48 sn103_48 202000.000000
Rwneg103_49 in103_49 sn103_49 202000.000000
Rwneg103_50 in103_50 sn103_50 78000.000000
Rwneg103_51 in103_51 sn103_51 202000.000000
Rwneg103_52 in103_52 sn103_52 202000.000000
Rwneg103_53 in103_53 sn103_53 78000.000000
Rwneg103_54 in103_54 sn103_54 202000.000000
Rwneg103_55 in103_55 sn103_55 202000.000000
Rwneg103_56 in103_56 sn103_56 202000.000000
Rwneg103_57 in103_57 sn103_57 202000.000000
Rwneg103_58 in103_58 sn103_58 78000.000000
Rwneg103_59 in103_59 sn103_59 78000.000000
Rwneg103_60 in103_60 sn103_60 78000.000000
Rwneg103_61 in103_61 sn103_61 78000.000000
Rwneg103_62 in103_62 sn103_62 202000.000000
Rwneg103_63 in103_63 sn103_63 202000.000000
Rwneg103_64 in103_64 sn103_64 202000.000000
Rwneg103_65 in103_65 sn103_65 78000.000000
Rwneg103_66 in103_66 sn103_66 78000.000000
Rwneg103_67 in103_67 sn103_67 78000.000000
Rwneg103_68 in103_68 sn103_68 78000.000000
Rwneg103_69 in103_69 sn103_69 202000.000000
Rwneg103_70 in103_70 sn103_70 202000.000000
Rwneg103_71 in103_71 sn103_71 202000.000000
Rwneg103_72 in103_72 sn103_72 202000.000000
Rwneg103_73 in103_73 sn103_73 202000.000000
Rwneg103_74 in103_74 sn103_74 78000.000000
Rwneg103_75 in103_75 sn103_75 202000.000000
Rwneg103_76 in103_76 sn103_76 202000.000000
Rwneg103_77 in103_77 sn103_77 202000.000000
Rwneg103_78 in103_78 sn103_78 78000.000000
Rwneg103_79 in103_79 sn103_79 202000.000000
Rwneg103_80 in103_80 sn103_80 202000.000000
Rwneg103_81 in103_81 sn103_81 202000.000000
Rwneg103_82 in103_82 sn103_82 78000.000000
Rwneg103_83 in103_83 sn103_83 78000.000000
Rwneg103_84 in103_84 sn103_84 202000.000000
Rwneg104_1 in104_1 sn104_1 202000.000000
Rwneg104_2 in104_2 sn104_2 202000.000000
Rwneg104_3 in104_3 sn104_3 202000.000000
Rwneg104_4 in104_4 sn104_4 202000.000000
Rwneg104_5 in104_5 sn104_5 78000.000000
Rwneg104_6 in104_6 sn104_6 78000.000000
Rwneg104_7 in104_7 sn104_7 202000.000000
Rwneg104_8 in104_8 sn104_8 202000.000000
Rwneg104_9 in104_9 sn104_9 78000.000000
Rwneg104_10 in104_10 sn104_10 78000.000000
Rwneg104_11 in104_11 sn104_11 202000.000000
Rwneg104_12 in104_12 sn104_12 78000.000000
Rwneg104_13 in104_13 sn104_13 78000.000000
Rwneg104_14 in104_14 sn104_14 202000.000000
Rwneg104_15 in104_15 sn104_15 202000.000000
Rwneg104_16 in104_16 sn104_16 202000.000000
Rwneg104_17 in104_17 sn104_17 78000.000000
Rwneg104_18 in104_18 sn104_18 78000.000000
Rwneg104_19 in104_19 sn104_19 202000.000000
Rwneg104_20 in104_20 sn104_20 202000.000000
Rwneg104_21 in104_21 sn104_21 78000.000000
Rwneg104_22 in104_22 sn104_22 202000.000000
Rwneg104_23 in104_23 sn104_23 202000.000000
Rwneg104_24 in104_24 sn104_24 78000.000000
Rwneg104_25 in104_25 sn104_25 202000.000000
Rwneg104_26 in104_26 sn104_26 78000.000000
Rwneg104_27 in104_27 sn104_27 78000.000000
Rwneg104_28 in104_28 sn104_28 78000.000000
Rwneg104_29 in104_29 sn104_29 202000.000000
Rwneg104_30 in104_30 sn104_30 202000.000000
Rwneg104_31 in104_31 sn104_31 78000.000000
Rwneg104_32 in104_32 sn104_32 202000.000000
Rwneg104_33 in104_33 sn104_33 202000.000000
Rwneg104_34 in104_34 sn104_34 202000.000000
Rwneg104_35 in104_35 sn104_35 202000.000000
Rwneg104_36 in104_36 sn104_36 78000.000000
Rwneg104_37 in104_37 sn104_37 202000.000000
Rwneg104_38 in104_38 sn104_38 202000.000000
Rwneg104_39 in104_39 sn104_39 78000.000000
Rwneg104_40 in104_40 sn104_40 202000.000000
Rwneg104_41 in104_41 sn104_41 78000.000000
Rwneg104_42 in104_42 sn104_42 202000.000000
Rwneg104_43 in104_43 sn104_43 78000.000000
Rwneg104_44 in104_44 sn104_44 78000.000000
Rwneg104_45 in104_45 sn104_45 202000.000000
Rwneg104_46 in104_46 sn104_46 202000.000000
Rwneg104_47 in104_47 sn104_47 78000.000000
Rwneg104_48 in104_48 sn104_48 78000.000000
Rwneg104_49 in104_49 sn104_49 202000.000000
Rwneg104_50 in104_50 sn104_50 202000.000000
Rwneg104_51 in104_51 sn104_51 78000.000000
Rwneg104_52 in104_52 sn104_52 202000.000000
Rwneg104_53 in104_53 sn104_53 202000.000000
Rwneg104_54 in104_54 sn104_54 78000.000000
Rwneg104_55 in104_55 sn104_55 202000.000000
Rwneg104_56 in104_56 sn104_56 78000.000000
Rwneg104_57 in104_57 sn104_57 202000.000000
Rwneg104_58 in104_58 sn104_58 202000.000000
Rwneg104_59 in104_59 sn104_59 202000.000000
Rwneg104_60 in104_60 sn104_60 78000.000000
Rwneg104_61 in104_61 sn104_61 202000.000000
Rwneg104_62 in104_62 sn104_62 78000.000000
Rwneg104_63 in104_63 sn104_63 78000.000000
Rwneg104_64 in104_64 sn104_64 78000.000000
Rwneg104_65 in104_65 sn104_65 78000.000000
Rwneg104_66 in104_66 sn104_66 202000.000000
Rwneg104_67 in104_67 sn104_67 78000.000000
Rwneg104_68 in104_68 sn104_68 78000.000000
Rwneg104_69 in104_69 sn104_69 78000.000000
Rwneg104_70 in104_70 sn104_70 202000.000000
Rwneg104_71 in104_71 sn104_71 202000.000000
Rwneg104_72 in104_72 sn104_72 78000.000000
Rwneg104_73 in104_73 sn104_73 202000.000000
Rwneg104_74 in104_74 sn104_74 202000.000000
Rwneg104_75 in104_75 sn104_75 202000.000000
Rwneg104_76 in104_76 sn104_76 202000.000000
Rwneg104_77 in104_77 sn104_77 78000.000000
Rwneg104_78 in104_78 sn104_78 78000.000000
Rwneg104_79 in104_79 sn104_79 78000.000000
Rwneg104_80 in104_80 sn104_80 78000.000000
Rwneg104_81 in104_81 sn104_81 78000.000000
Rwneg104_82 in104_82 sn104_82 78000.000000
Rwneg104_83 in104_83 sn104_83 202000.000000
Rwneg104_84 in104_84 sn104_84 202000.000000
Rwneg105_1 in105_1 sn105_1 78000.000000
Rwneg105_2 in105_2 sn105_2 202000.000000
Rwneg105_3 in105_3 sn105_3 202000.000000
Rwneg105_4 in105_4 sn105_4 202000.000000
Rwneg105_5 in105_5 sn105_5 202000.000000
Rwneg105_6 in105_6 sn105_6 78000.000000
Rwneg105_7 in105_7 sn105_7 78000.000000
Rwneg105_8 in105_8 sn105_8 202000.000000
Rwneg105_9 in105_9 sn105_9 202000.000000
Rwneg105_10 in105_10 sn105_10 202000.000000
Rwneg105_11 in105_11 sn105_11 78000.000000
Rwneg105_12 in105_12 sn105_12 202000.000000
Rwneg105_13 in105_13 sn105_13 78000.000000
Rwneg105_14 in105_14 sn105_14 78000.000000
Rwneg105_15 in105_15 sn105_15 78000.000000
Rwneg105_16 in105_16 sn105_16 202000.000000
Rwneg105_17 in105_17 sn105_17 78000.000000
Rwneg105_18 in105_18 sn105_18 202000.000000
Rwneg105_19 in105_19 sn105_19 202000.000000
Rwneg105_20 in105_20 sn105_20 202000.000000
Rwneg105_21 in105_21 sn105_21 78000.000000
Rwneg105_22 in105_22 sn105_22 78000.000000
Rwneg105_23 in105_23 sn105_23 78000.000000
Rwneg105_24 in105_24 sn105_24 78000.000000
Rwneg105_25 in105_25 sn105_25 202000.000000
Rwneg105_26 in105_26 sn105_26 78000.000000
Rwneg105_27 in105_27 sn105_27 202000.000000
Rwneg105_28 in105_28 sn105_28 78000.000000
Rwneg105_29 in105_29 sn105_29 202000.000000
Rwneg105_30 in105_30 sn105_30 78000.000000
Rwneg105_31 in105_31 sn105_31 78000.000000
Rwneg105_32 in105_32 sn105_32 202000.000000
Rwneg105_33 in105_33 sn105_33 78000.000000
Rwneg105_34 in105_34 sn105_34 202000.000000
Rwneg105_35 in105_35 sn105_35 202000.000000
Rwneg105_36 in105_36 sn105_36 202000.000000
Rwneg105_37 in105_37 sn105_37 202000.000000
Rwneg105_38 in105_38 sn105_38 202000.000000
Rwneg105_39 in105_39 sn105_39 202000.000000
Rwneg105_40 in105_40 sn105_40 202000.000000
Rwneg105_41 in105_41 sn105_41 78000.000000
Rwneg105_42 in105_42 sn105_42 202000.000000
Rwneg105_43 in105_43 sn105_43 78000.000000
Rwneg105_44 in105_44 sn105_44 78000.000000
Rwneg105_45 in105_45 sn105_45 202000.000000
Rwneg105_46 in105_46 sn105_46 78000.000000
Rwneg105_47 in105_47 sn105_47 78000.000000
Rwneg105_48 in105_48 sn105_48 78000.000000
Rwneg105_49 in105_49 sn105_49 202000.000000
Rwneg105_50 in105_50 sn105_50 202000.000000
Rwneg105_51 in105_51 sn105_51 202000.000000
Rwneg105_52 in105_52 sn105_52 202000.000000
Rwneg105_53 in105_53 sn105_53 202000.000000
Rwneg105_54 in105_54 sn105_54 202000.000000
Rwneg105_55 in105_55 sn105_55 202000.000000
Rwneg105_56 in105_56 sn105_56 202000.000000
Rwneg105_57 in105_57 sn105_57 78000.000000
Rwneg105_58 in105_58 sn105_58 202000.000000
Rwneg105_59 in105_59 sn105_59 202000.000000
Rwneg105_60 in105_60 sn105_60 78000.000000
Rwneg105_61 in105_61 sn105_61 202000.000000
Rwneg105_62 in105_62 sn105_62 78000.000000
Rwneg105_63 in105_63 sn105_63 202000.000000
Rwneg105_64 in105_64 sn105_64 202000.000000
Rwneg105_65 in105_65 sn105_65 202000.000000
Rwneg105_66 in105_66 sn105_66 202000.000000
Rwneg105_67 in105_67 sn105_67 202000.000000
Rwneg105_68 in105_68 sn105_68 78000.000000
Rwneg105_69 in105_69 sn105_69 202000.000000
Rwneg105_70 in105_70 sn105_70 202000.000000
Rwneg105_71 in105_71 sn105_71 202000.000000
Rwneg105_72 in105_72 sn105_72 78000.000000
Rwneg105_73 in105_73 sn105_73 78000.000000
Rwneg105_74 in105_74 sn105_74 202000.000000
Rwneg105_75 in105_75 sn105_75 202000.000000
Rwneg105_76 in105_76 sn105_76 202000.000000
Rwneg105_77 in105_77 sn105_77 202000.000000
Rwneg105_78 in105_78 sn105_78 78000.000000
Rwneg105_79 in105_79 sn105_79 202000.000000
Rwneg105_80 in105_80 sn105_80 202000.000000
Rwneg105_81 in105_81 sn105_81 78000.000000
Rwneg105_82 in105_82 sn105_82 202000.000000
Rwneg105_83 in105_83 sn105_83 202000.000000
Rwneg105_84 in105_84 sn105_84 202000.000000
Rwneg106_1 in106_1 sn106_1 202000.000000
Rwneg106_2 in106_2 sn106_2 202000.000000
Rwneg106_3 in106_3 sn106_3 78000.000000
Rwneg106_4 in106_4 sn106_4 202000.000000
Rwneg106_5 in106_5 sn106_5 78000.000000
Rwneg106_6 in106_6 sn106_6 202000.000000
Rwneg106_7 in106_7 sn106_7 202000.000000
Rwneg106_8 in106_8 sn106_8 78000.000000
Rwneg106_9 in106_9 sn106_9 78000.000000
Rwneg106_10 in106_10 sn106_10 202000.000000
Rwneg106_11 in106_11 sn106_11 78000.000000
Rwneg106_12 in106_12 sn106_12 202000.000000
Rwneg106_13 in106_13 sn106_13 78000.000000
Rwneg106_14 in106_14 sn106_14 202000.000000
Rwneg106_15 in106_15 sn106_15 78000.000000
Rwneg106_16 in106_16 sn106_16 202000.000000
Rwneg106_17 in106_17 sn106_17 202000.000000
Rwneg106_18 in106_18 sn106_18 78000.000000
Rwneg106_19 in106_19 sn106_19 202000.000000
Rwneg106_20 in106_20 sn106_20 78000.000000
Rwneg106_21 in106_21 sn106_21 78000.000000
Rwneg106_22 in106_22 sn106_22 202000.000000
Rwneg106_23 in106_23 sn106_23 78000.000000
Rwneg106_24 in106_24 sn106_24 202000.000000
Rwneg106_25 in106_25 sn106_25 78000.000000
Rwneg106_26 in106_26 sn106_26 78000.000000
Rwneg106_27 in106_27 sn106_27 202000.000000
Rwneg106_28 in106_28 sn106_28 202000.000000
Rwneg106_29 in106_29 sn106_29 78000.000000
Rwneg106_30 in106_30 sn106_30 202000.000000
Rwneg106_31 in106_31 sn106_31 202000.000000
Rwneg106_32 in106_32 sn106_32 202000.000000
Rwneg106_33 in106_33 sn106_33 78000.000000
Rwneg106_34 in106_34 sn106_34 78000.000000
Rwneg106_35 in106_35 sn106_35 78000.000000
Rwneg106_36 in106_36 sn106_36 202000.000000
Rwneg106_37 in106_37 sn106_37 202000.000000
Rwneg106_38 in106_38 sn106_38 202000.000000
Rwneg106_39 in106_39 sn106_39 78000.000000
Rwneg106_40 in106_40 sn106_40 202000.000000
Rwneg106_41 in106_41 sn106_41 78000.000000
Rwneg106_42 in106_42 sn106_42 202000.000000
Rwneg106_43 in106_43 sn106_43 78000.000000
Rwneg106_44 in106_44 sn106_44 202000.000000
Rwneg106_45 in106_45 sn106_45 202000.000000
Rwneg106_46 in106_46 sn106_46 202000.000000
Rwneg106_47 in106_47 sn106_47 202000.000000
Rwneg106_48 in106_48 sn106_48 78000.000000
Rwneg106_49 in106_49 sn106_49 202000.000000
Rwneg106_50 in106_50 sn106_50 202000.000000
Rwneg106_51 in106_51 sn106_51 202000.000000
Rwneg106_52 in106_52 sn106_52 202000.000000
Rwneg106_53 in106_53 sn106_53 78000.000000
Rwneg106_54 in106_54 sn106_54 202000.000000
Rwneg106_55 in106_55 sn106_55 78000.000000
Rwneg106_56 in106_56 sn106_56 78000.000000
Rwneg106_57 in106_57 sn106_57 202000.000000
Rwneg106_58 in106_58 sn106_58 202000.000000
Rwneg106_59 in106_59 sn106_59 78000.000000
Rwneg106_60 in106_60 sn106_60 202000.000000
Rwneg106_61 in106_61 sn106_61 78000.000000
Rwneg106_62 in106_62 sn106_62 202000.000000
Rwneg106_63 in106_63 sn106_63 78000.000000
Rwneg106_64 in106_64 sn106_64 78000.000000
Rwneg106_65 in106_65 sn106_65 78000.000000
Rwneg106_66 in106_66 sn106_66 202000.000000
Rwneg106_67 in106_67 sn106_67 202000.000000
Rwneg106_68 in106_68 sn106_68 202000.000000
Rwneg106_69 in106_69 sn106_69 78000.000000
Rwneg106_70 in106_70 sn106_70 202000.000000
Rwneg106_71 in106_71 sn106_71 78000.000000
Rwneg106_72 in106_72 sn106_72 202000.000000
Rwneg106_73 in106_73 sn106_73 78000.000000
Rwneg106_74 in106_74 sn106_74 78000.000000
Rwneg106_75 in106_75 sn106_75 78000.000000
Rwneg106_76 in106_76 sn106_76 202000.000000
Rwneg106_77 in106_77 sn106_77 78000.000000
Rwneg106_78 in106_78 sn106_78 202000.000000
Rwneg106_79 in106_79 sn106_79 78000.000000
Rwneg106_80 in106_80 sn106_80 78000.000000
Rwneg106_81 in106_81 sn106_81 78000.000000
Rwneg106_82 in106_82 sn106_82 78000.000000
Rwneg106_83 in106_83 sn106_83 78000.000000
Rwneg106_84 in106_84 sn106_84 78000.000000
Rwneg107_1 in107_1 sn107_1 202000.000000
Rwneg107_2 in107_2 sn107_2 202000.000000
Rwneg107_3 in107_3 sn107_3 202000.000000
Rwneg107_4 in107_4 sn107_4 202000.000000
Rwneg107_5 in107_5 sn107_5 202000.000000
Rwneg107_6 in107_6 sn107_6 202000.000000
Rwneg107_7 in107_7 sn107_7 78000.000000
Rwneg107_8 in107_8 sn107_8 78000.000000
Rwneg107_9 in107_9 sn107_9 202000.000000
Rwneg107_10 in107_10 sn107_10 78000.000000
Rwneg107_11 in107_11 sn107_11 78000.000000
Rwneg107_12 in107_12 sn107_12 78000.000000
Rwneg107_13 in107_13 sn107_13 202000.000000
Rwneg107_14 in107_14 sn107_14 202000.000000
Rwneg107_15 in107_15 sn107_15 202000.000000
Rwneg107_16 in107_16 sn107_16 202000.000000
Rwneg107_17 in107_17 sn107_17 202000.000000
Rwneg107_18 in107_18 sn107_18 78000.000000
Rwneg107_19 in107_19 sn107_19 202000.000000
Rwneg107_20 in107_20 sn107_20 78000.000000
Rwneg107_21 in107_21 sn107_21 202000.000000
Rwneg107_22 in107_22 sn107_22 202000.000000
Rwneg107_23 in107_23 sn107_23 78000.000000
Rwneg107_24 in107_24 sn107_24 202000.000000
Rwneg107_25 in107_25 sn107_25 202000.000000
Rwneg107_26 in107_26 sn107_26 202000.000000
Rwneg107_27 in107_27 sn107_27 202000.000000
Rwneg107_28 in107_28 sn107_28 202000.000000
Rwneg107_29 in107_29 sn107_29 78000.000000
Rwneg107_30 in107_30 sn107_30 202000.000000
Rwneg107_31 in107_31 sn107_31 202000.000000
Rwneg107_32 in107_32 sn107_32 78000.000000
Rwneg107_33 in107_33 sn107_33 202000.000000
Rwneg107_34 in107_34 sn107_34 78000.000000
Rwneg107_35 in107_35 sn107_35 202000.000000
Rwneg107_36 in107_36 sn107_36 78000.000000
Rwneg107_37 in107_37 sn107_37 78000.000000
Rwneg107_38 in107_38 sn107_38 202000.000000
Rwneg107_39 in107_39 sn107_39 78000.000000
Rwneg107_40 in107_40 sn107_40 78000.000000
Rwneg107_41 in107_41 sn107_41 202000.000000
Rwneg107_42 in107_42 sn107_42 202000.000000
Rwneg107_43 in107_43 sn107_43 202000.000000
Rwneg107_44 in107_44 sn107_44 202000.000000
Rwneg107_45 in107_45 sn107_45 202000.000000
Rwneg107_46 in107_46 sn107_46 78000.000000
Rwneg107_47 in107_47 sn107_47 202000.000000
Rwneg107_48 in107_48 sn107_48 78000.000000
Rwneg107_49 in107_49 sn107_49 78000.000000
Rwneg107_50 in107_50 sn107_50 202000.000000
Rwneg107_51 in107_51 sn107_51 202000.000000
Rwneg107_52 in107_52 sn107_52 78000.000000
Rwneg107_53 in107_53 sn107_53 78000.000000
Rwneg107_54 in107_54 sn107_54 202000.000000
Rwneg107_55 in107_55 sn107_55 78000.000000
Rwneg107_56 in107_56 sn107_56 78000.000000
Rwneg107_57 in107_57 sn107_57 78000.000000
Rwneg107_58 in107_58 sn107_58 78000.000000
Rwneg107_59 in107_59 sn107_59 202000.000000
Rwneg107_60 in107_60 sn107_60 202000.000000
Rwneg107_61 in107_61 sn107_61 78000.000000
Rwneg107_62 in107_62 sn107_62 202000.000000
Rwneg107_63 in107_63 sn107_63 78000.000000
Rwneg107_64 in107_64 sn107_64 78000.000000
Rwneg107_65 in107_65 sn107_65 78000.000000
Rwneg107_66 in107_66 sn107_66 78000.000000
Rwneg107_67 in107_67 sn107_67 202000.000000
Rwneg107_68 in107_68 sn107_68 78000.000000
Rwneg107_69 in107_69 sn107_69 78000.000000
Rwneg107_70 in107_70 sn107_70 202000.000000
Rwneg107_71 in107_71 sn107_71 78000.000000
Rwneg107_72 in107_72 sn107_72 202000.000000
Rwneg107_73 in107_73 sn107_73 78000.000000
Rwneg107_74 in107_74 sn107_74 202000.000000
Rwneg107_75 in107_75 sn107_75 78000.000000
Rwneg107_76 in107_76 sn107_76 78000.000000
Rwneg107_77 in107_77 sn107_77 78000.000000
Rwneg107_78 in107_78 sn107_78 202000.000000
Rwneg107_79 in107_79 sn107_79 78000.000000
Rwneg107_80 in107_80 sn107_80 78000.000000
Rwneg107_81 in107_81 sn107_81 202000.000000
Rwneg107_82 in107_82 sn107_82 78000.000000
Rwneg107_83 in107_83 sn107_83 78000.000000
Rwneg107_84 in107_84 sn107_84 202000.000000
Rwneg108_1 in108_1 sn108_1 202000.000000
Rwneg108_2 in108_2 sn108_2 202000.000000
Rwneg108_3 in108_3 sn108_3 202000.000000
Rwneg108_4 in108_4 sn108_4 202000.000000
Rwneg108_5 in108_5 sn108_5 202000.000000
Rwneg108_6 in108_6 sn108_6 202000.000000
Rwneg108_7 in108_7 sn108_7 202000.000000
Rwneg108_8 in108_8 sn108_8 202000.000000
Rwneg108_9 in108_9 sn108_9 202000.000000
Rwneg108_10 in108_10 sn108_10 78000.000000
Rwneg108_11 in108_11 sn108_11 202000.000000
Rwneg108_12 in108_12 sn108_12 202000.000000
Rwneg108_13 in108_13 sn108_13 202000.000000
Rwneg108_14 in108_14 sn108_14 202000.000000
Rwneg108_15 in108_15 sn108_15 78000.000000
Rwneg108_16 in108_16 sn108_16 78000.000000
Rwneg108_17 in108_17 sn108_17 202000.000000
Rwneg108_18 in108_18 sn108_18 78000.000000
Rwneg108_19 in108_19 sn108_19 78000.000000
Rwneg108_20 in108_20 sn108_20 78000.000000
Rwneg108_21 in108_21 sn108_21 202000.000000
Rwneg108_22 in108_22 sn108_22 202000.000000
Rwneg108_23 in108_23 sn108_23 78000.000000
Rwneg108_24 in108_24 sn108_24 202000.000000
Rwneg108_25 in108_25 sn108_25 78000.000000
Rwneg108_26 in108_26 sn108_26 78000.000000
Rwneg108_27 in108_27 sn108_27 202000.000000
Rwneg108_28 in108_28 sn108_28 78000.000000
Rwneg108_29 in108_29 sn108_29 202000.000000
Rwneg108_30 in108_30 sn108_30 202000.000000
Rwneg108_31 in108_31 sn108_31 202000.000000
Rwneg108_32 in108_32 sn108_32 202000.000000
Rwneg108_33 in108_33 sn108_33 78000.000000
Rwneg108_34 in108_34 sn108_34 202000.000000
Rwneg108_35 in108_35 sn108_35 202000.000000
Rwneg108_36 in108_36 sn108_36 202000.000000
Rwneg108_37 in108_37 sn108_37 78000.000000
Rwneg108_38 in108_38 sn108_38 78000.000000
Rwneg108_39 in108_39 sn108_39 78000.000000
Rwneg108_40 in108_40 sn108_40 78000.000000
Rwneg108_41 in108_41 sn108_41 78000.000000
Rwneg108_42 in108_42 sn108_42 202000.000000
Rwneg108_43 in108_43 sn108_43 78000.000000
Rwneg108_44 in108_44 sn108_44 202000.000000
Rwneg108_45 in108_45 sn108_45 78000.000000
Rwneg108_46 in108_46 sn108_46 202000.000000
Rwneg108_47 in108_47 sn108_47 202000.000000
Rwneg108_48 in108_48 sn108_48 202000.000000
Rwneg108_49 in108_49 sn108_49 78000.000000
Rwneg108_50 in108_50 sn108_50 202000.000000
Rwneg108_51 in108_51 sn108_51 78000.000000
Rwneg108_52 in108_52 sn108_52 202000.000000
Rwneg108_53 in108_53 sn108_53 78000.000000
Rwneg108_54 in108_54 sn108_54 202000.000000
Rwneg108_55 in108_55 sn108_55 78000.000000
Rwneg108_56 in108_56 sn108_56 78000.000000
Rwneg108_57 in108_57 sn108_57 202000.000000
Rwneg108_58 in108_58 sn108_58 202000.000000
Rwneg108_59 in108_59 sn108_59 202000.000000
Rwneg108_60 in108_60 sn108_60 202000.000000
Rwneg108_61 in108_61 sn108_61 202000.000000
Rwneg108_62 in108_62 sn108_62 202000.000000
Rwneg108_63 in108_63 sn108_63 78000.000000
Rwneg108_64 in108_64 sn108_64 78000.000000
Rwneg108_65 in108_65 sn108_65 78000.000000
Rwneg108_66 in108_66 sn108_66 202000.000000
Rwneg108_67 in108_67 sn108_67 202000.000000
Rwneg108_68 in108_68 sn108_68 202000.000000
Rwneg108_69 in108_69 sn108_69 202000.000000
Rwneg108_70 in108_70 sn108_70 78000.000000
Rwneg108_71 in108_71 sn108_71 78000.000000
Rwneg108_72 in108_72 sn108_72 202000.000000
Rwneg108_73 in108_73 sn108_73 202000.000000
Rwneg108_74 in108_74 sn108_74 202000.000000
Rwneg108_75 in108_75 sn108_75 78000.000000
Rwneg108_76 in108_76 sn108_76 202000.000000
Rwneg108_77 in108_77 sn108_77 78000.000000
Rwneg108_78 in108_78 sn108_78 202000.000000
Rwneg108_79 in108_79 sn108_79 202000.000000
Rwneg108_80 in108_80 sn108_80 78000.000000
Rwneg108_81 in108_81 sn108_81 202000.000000
Rwneg108_82 in108_82 sn108_82 202000.000000
Rwneg108_83 in108_83 sn108_83 202000.000000
Rwneg108_84 in108_84 sn108_84 78000.000000
Rwneg109_1 in109_1 sn109_1 78000.000000
Rwneg109_2 in109_2 sn109_2 78000.000000
Rwneg109_3 in109_3 sn109_3 78000.000000
Rwneg109_4 in109_4 sn109_4 78000.000000
Rwneg109_5 in109_5 sn109_5 78000.000000
Rwneg109_6 in109_6 sn109_6 78000.000000
Rwneg109_7 in109_7 sn109_7 202000.000000
Rwneg109_8 in109_8 sn109_8 78000.000000
Rwneg109_9 in109_9 sn109_9 202000.000000
Rwneg109_10 in109_10 sn109_10 202000.000000
Rwneg109_11 in109_11 sn109_11 202000.000000
Rwneg109_12 in109_12 sn109_12 78000.000000
Rwneg109_13 in109_13 sn109_13 78000.000000
Rwneg109_14 in109_14 sn109_14 78000.000000
Rwneg109_15 in109_15 sn109_15 202000.000000
Rwneg109_16 in109_16 sn109_16 78000.000000
Rwneg109_17 in109_17 sn109_17 202000.000000
Rwneg109_18 in109_18 sn109_18 78000.000000
Rwneg109_19 in109_19 sn109_19 78000.000000
Rwneg109_20 in109_20 sn109_20 202000.000000
Rwneg109_21 in109_21 sn109_21 78000.000000
Rwneg109_22 in109_22 sn109_22 78000.000000
Rwneg109_23 in109_23 sn109_23 202000.000000
Rwneg109_24 in109_24 sn109_24 202000.000000
Rwneg109_25 in109_25 sn109_25 78000.000000
Rwneg109_26 in109_26 sn109_26 202000.000000
Rwneg109_27 in109_27 sn109_27 78000.000000
Rwneg109_28 in109_28 sn109_28 202000.000000
Rwneg109_29 in109_29 sn109_29 202000.000000
Rwneg109_30 in109_30 sn109_30 78000.000000
Rwneg109_31 in109_31 sn109_31 78000.000000
Rwneg109_32 in109_32 sn109_32 202000.000000
Rwneg109_33 in109_33 sn109_33 202000.000000
Rwneg109_34 in109_34 sn109_34 202000.000000
Rwneg109_35 in109_35 sn109_35 78000.000000
Rwneg109_36 in109_36 sn109_36 202000.000000
Rwneg109_37 in109_37 sn109_37 202000.000000
Rwneg109_38 in109_38 sn109_38 78000.000000
Rwneg109_39 in109_39 sn109_39 78000.000000
Rwneg109_40 in109_40 sn109_40 202000.000000
Rwneg109_41 in109_41 sn109_41 78000.000000
Rwneg109_42 in109_42 sn109_42 78000.000000
Rwneg109_43 in109_43 sn109_43 78000.000000
Rwneg109_44 in109_44 sn109_44 78000.000000
Rwneg109_45 in109_45 sn109_45 78000.000000
Rwneg109_46 in109_46 sn109_46 202000.000000
Rwneg109_47 in109_47 sn109_47 78000.000000
Rwneg109_48 in109_48 sn109_48 78000.000000
Rwneg109_49 in109_49 sn109_49 78000.000000
Rwneg109_50 in109_50 sn109_50 202000.000000
Rwneg109_51 in109_51 sn109_51 202000.000000
Rwneg109_52 in109_52 sn109_52 202000.000000
Rwneg109_53 in109_53 sn109_53 202000.000000
Rwneg109_54 in109_54 sn109_54 202000.000000
Rwneg109_55 in109_55 sn109_55 78000.000000
Rwneg109_56 in109_56 sn109_56 202000.000000
Rwneg109_57 in109_57 sn109_57 202000.000000
Rwneg109_58 in109_58 sn109_58 202000.000000
Rwneg109_59 in109_59 sn109_59 78000.000000
Rwneg109_60 in109_60 sn109_60 202000.000000
Rwneg109_61 in109_61 sn109_61 78000.000000
Rwneg109_62 in109_62 sn109_62 202000.000000
Rwneg109_63 in109_63 sn109_63 202000.000000
Rwneg109_64 in109_64 sn109_64 78000.000000
Rwneg109_65 in109_65 sn109_65 202000.000000
Rwneg109_66 in109_66 sn109_66 202000.000000
Rwneg109_67 in109_67 sn109_67 78000.000000
Rwneg109_68 in109_68 sn109_68 202000.000000
Rwneg109_69 in109_69 sn109_69 202000.000000
Rwneg109_70 in109_70 sn109_70 78000.000000
Rwneg109_71 in109_71 sn109_71 202000.000000
Rwneg109_72 in109_72 sn109_72 78000.000000
Rwneg109_73 in109_73 sn109_73 202000.000000
Rwneg109_74 in109_74 sn109_74 78000.000000
Rwneg109_75 in109_75 sn109_75 78000.000000
Rwneg109_76 in109_76 sn109_76 78000.000000
Rwneg109_77 in109_77 sn109_77 202000.000000
Rwneg109_78 in109_78 sn109_78 202000.000000
Rwneg109_79 in109_79 sn109_79 202000.000000
Rwneg109_80 in109_80 sn109_80 202000.000000
Rwneg109_81 in109_81 sn109_81 202000.000000
Rwneg109_82 in109_82 sn109_82 202000.000000
Rwneg109_83 in109_83 sn109_83 78000.000000
Rwneg109_84 in109_84 sn109_84 202000.000000
Rwneg110_1 in110_1 sn110_1 202000.000000
Rwneg110_2 in110_2 sn110_2 78000.000000
Rwneg110_3 in110_3 sn110_3 202000.000000
Rwneg110_4 in110_4 sn110_4 202000.000000
Rwneg110_5 in110_5 sn110_5 202000.000000
Rwneg110_6 in110_6 sn110_6 78000.000000
Rwneg110_7 in110_7 sn110_7 78000.000000
Rwneg110_8 in110_8 sn110_8 78000.000000
Rwneg110_9 in110_9 sn110_9 202000.000000
Rwneg110_10 in110_10 sn110_10 202000.000000
Rwneg110_11 in110_11 sn110_11 202000.000000
Rwneg110_12 in110_12 sn110_12 78000.000000
Rwneg110_13 in110_13 sn110_13 202000.000000
Rwneg110_14 in110_14 sn110_14 78000.000000
Rwneg110_15 in110_15 sn110_15 78000.000000
Rwneg110_16 in110_16 sn110_16 78000.000000
Rwneg110_17 in110_17 sn110_17 202000.000000
Rwneg110_18 in110_18 sn110_18 202000.000000
Rwneg110_19 in110_19 sn110_19 78000.000000
Rwneg110_20 in110_20 sn110_20 78000.000000
Rwneg110_21 in110_21 sn110_21 202000.000000
Rwneg110_22 in110_22 sn110_22 202000.000000
Rwneg110_23 in110_23 sn110_23 202000.000000
Rwneg110_24 in110_24 sn110_24 202000.000000
Rwneg110_25 in110_25 sn110_25 78000.000000
Rwneg110_26 in110_26 sn110_26 202000.000000
Rwneg110_27 in110_27 sn110_27 78000.000000
Rwneg110_28 in110_28 sn110_28 78000.000000
Rwneg110_29 in110_29 sn110_29 78000.000000
Rwneg110_30 in110_30 sn110_30 202000.000000
Rwneg110_31 in110_31 sn110_31 202000.000000
Rwneg110_32 in110_32 sn110_32 78000.000000
Rwneg110_33 in110_33 sn110_33 202000.000000
Rwneg110_34 in110_34 sn110_34 78000.000000
Rwneg110_35 in110_35 sn110_35 202000.000000
Rwneg110_36 in110_36 sn110_36 78000.000000
Rwneg110_37 in110_37 sn110_37 78000.000000
Rwneg110_38 in110_38 sn110_38 78000.000000
Rwneg110_39 in110_39 sn110_39 78000.000000
Rwneg110_40 in110_40 sn110_40 78000.000000
Rwneg110_41 in110_41 sn110_41 78000.000000
Rwneg110_42 in110_42 sn110_42 78000.000000
Rwneg110_43 in110_43 sn110_43 202000.000000
Rwneg110_44 in110_44 sn110_44 202000.000000
Rwneg110_45 in110_45 sn110_45 78000.000000
Rwneg110_46 in110_46 sn110_46 78000.000000
Rwneg110_47 in110_47 sn110_47 202000.000000
Rwneg110_48 in110_48 sn110_48 202000.000000
Rwneg110_49 in110_49 sn110_49 78000.000000
Rwneg110_50 in110_50 sn110_50 78000.000000
Rwneg110_51 in110_51 sn110_51 78000.000000
Rwneg110_52 in110_52 sn110_52 78000.000000
Rwneg110_53 in110_53 sn110_53 202000.000000
Rwneg110_54 in110_54 sn110_54 202000.000000
Rwneg110_55 in110_55 sn110_55 202000.000000
Rwneg110_56 in110_56 sn110_56 202000.000000
Rwneg110_57 in110_57 sn110_57 202000.000000
Rwneg110_58 in110_58 sn110_58 202000.000000
Rwneg110_59 in110_59 sn110_59 202000.000000
Rwneg110_60 in110_60 sn110_60 202000.000000
Rwneg110_61 in110_61 sn110_61 202000.000000
Rwneg110_62 in110_62 sn110_62 202000.000000
Rwneg110_63 in110_63 sn110_63 78000.000000
Rwneg110_64 in110_64 sn110_64 78000.000000
Rwneg110_65 in110_65 sn110_65 202000.000000
Rwneg110_66 in110_66 sn110_66 202000.000000
Rwneg110_67 in110_67 sn110_67 78000.000000
Rwneg110_68 in110_68 sn110_68 78000.000000
Rwneg110_69 in110_69 sn110_69 78000.000000
Rwneg110_70 in110_70 sn110_70 202000.000000
Rwneg110_71 in110_71 sn110_71 202000.000000
Rwneg110_72 in110_72 sn110_72 202000.000000
Rwneg110_73 in110_73 sn110_73 202000.000000
Rwneg110_74 in110_74 sn110_74 78000.000000
Rwneg110_75 in110_75 sn110_75 202000.000000
Rwneg110_76 in110_76 sn110_76 78000.000000
Rwneg110_77 in110_77 sn110_77 202000.000000
Rwneg110_78 in110_78 sn110_78 202000.000000
Rwneg110_79 in110_79 sn110_79 78000.000000
Rwneg110_80 in110_80 sn110_80 202000.000000
Rwneg110_81 in110_81 sn110_81 202000.000000
Rwneg110_82 in110_82 sn110_82 202000.000000
Rwneg110_83 in110_83 sn110_83 202000.000000
Rwneg110_84 in110_84 sn110_84 202000.000000
Rwneg111_1 in111_1 sn111_1 202000.000000
Rwneg111_2 in111_2 sn111_2 202000.000000
Rwneg111_3 in111_3 sn111_3 202000.000000
Rwneg111_4 in111_4 sn111_4 78000.000000
Rwneg111_5 in111_5 sn111_5 78000.000000
Rwneg111_6 in111_6 sn111_6 78000.000000
Rwneg111_7 in111_7 sn111_7 202000.000000
Rwneg111_8 in111_8 sn111_8 202000.000000
Rwneg111_9 in111_9 sn111_9 78000.000000
Rwneg111_10 in111_10 sn111_10 78000.000000
Rwneg111_11 in111_11 sn111_11 202000.000000
Rwneg111_12 in111_12 sn111_12 78000.000000
Rwneg111_13 in111_13 sn111_13 78000.000000
Rwneg111_14 in111_14 sn111_14 202000.000000
Rwneg111_15 in111_15 sn111_15 78000.000000
Rwneg111_16 in111_16 sn111_16 78000.000000
Rwneg111_17 in111_17 sn111_17 202000.000000
Rwneg111_18 in111_18 sn111_18 78000.000000
Rwneg111_19 in111_19 sn111_19 78000.000000
Rwneg111_20 in111_20 sn111_20 78000.000000
Rwneg111_21 in111_21 sn111_21 78000.000000
Rwneg111_22 in111_22 sn111_22 78000.000000
Rwneg111_23 in111_23 sn111_23 202000.000000
Rwneg111_24 in111_24 sn111_24 78000.000000
Rwneg111_25 in111_25 sn111_25 202000.000000
Rwneg111_26 in111_26 sn111_26 78000.000000
Rwneg111_27 in111_27 sn111_27 78000.000000
Rwneg111_28 in111_28 sn111_28 78000.000000
Rwneg111_29 in111_29 sn111_29 78000.000000
Rwneg111_30 in111_30 sn111_30 202000.000000
Rwneg111_31 in111_31 sn111_31 202000.000000
Rwneg111_32 in111_32 sn111_32 202000.000000
Rwneg111_33 in111_33 sn111_33 78000.000000
Rwneg111_34 in111_34 sn111_34 202000.000000
Rwneg111_35 in111_35 sn111_35 78000.000000
Rwneg111_36 in111_36 sn111_36 78000.000000
Rwneg111_37 in111_37 sn111_37 202000.000000
Rwneg111_38 in111_38 sn111_38 78000.000000
Rwneg111_39 in111_39 sn111_39 78000.000000
Rwneg111_40 in111_40 sn111_40 78000.000000
Rwneg111_41 in111_41 sn111_41 78000.000000
Rwneg111_42 in111_42 sn111_42 202000.000000
Rwneg111_43 in111_43 sn111_43 202000.000000
Rwneg111_44 in111_44 sn111_44 78000.000000
Rwneg111_45 in111_45 sn111_45 78000.000000
Rwneg111_46 in111_46 sn111_46 202000.000000
Rwneg111_47 in111_47 sn111_47 78000.000000
Rwneg111_48 in111_48 sn111_48 202000.000000
Rwneg111_49 in111_49 sn111_49 202000.000000
Rwneg111_50 in111_50 sn111_50 202000.000000
Rwneg111_51 in111_51 sn111_51 202000.000000
Rwneg111_52 in111_52 sn111_52 202000.000000
Rwneg111_53 in111_53 sn111_53 78000.000000
Rwneg111_54 in111_54 sn111_54 78000.000000
Rwneg111_55 in111_55 sn111_55 78000.000000
Rwneg111_56 in111_56 sn111_56 202000.000000
Rwneg111_57 in111_57 sn111_57 202000.000000
Rwneg111_58 in111_58 sn111_58 202000.000000
Rwneg111_59 in111_59 sn111_59 202000.000000
Rwneg111_60 in111_60 sn111_60 78000.000000
Rwneg111_61 in111_61 sn111_61 202000.000000
Rwneg111_62 in111_62 sn111_62 202000.000000
Rwneg111_63 in111_63 sn111_63 78000.000000
Rwneg111_64 in111_64 sn111_64 78000.000000
Rwneg111_65 in111_65 sn111_65 202000.000000
Rwneg111_66 in111_66 sn111_66 202000.000000
Rwneg111_67 in111_67 sn111_67 78000.000000
Rwneg111_68 in111_68 sn111_68 78000.000000
Rwneg111_69 in111_69 sn111_69 202000.000000
Rwneg111_70 in111_70 sn111_70 78000.000000
Rwneg111_71 in111_71 sn111_71 78000.000000
Rwneg111_72 in111_72 sn111_72 78000.000000
Rwneg111_73 in111_73 sn111_73 202000.000000
Rwneg111_74 in111_74 sn111_74 202000.000000
Rwneg111_75 in111_75 sn111_75 78000.000000
Rwneg111_76 in111_76 sn111_76 202000.000000
Rwneg111_77 in111_77 sn111_77 78000.000000
Rwneg111_78 in111_78 sn111_78 78000.000000
Rwneg111_79 in111_79 sn111_79 202000.000000
Rwneg111_80 in111_80 sn111_80 78000.000000
Rwneg111_81 in111_81 sn111_81 202000.000000
Rwneg111_82 in111_82 sn111_82 78000.000000
Rwneg111_83 in111_83 sn111_83 78000.000000
Rwneg111_84 in111_84 sn111_84 202000.000000
Rwneg112_1 in112_1 sn112_1 78000.000000
Rwneg112_2 in112_2 sn112_2 202000.000000
Rwneg112_3 in112_3 sn112_3 78000.000000
Rwneg112_4 in112_4 sn112_4 202000.000000
Rwneg112_5 in112_5 sn112_5 78000.000000
Rwneg112_6 in112_6 sn112_6 78000.000000
Rwneg112_7 in112_7 sn112_7 202000.000000
Rwneg112_8 in112_8 sn112_8 78000.000000
Rwneg112_9 in112_9 sn112_9 78000.000000
Rwneg112_10 in112_10 sn112_10 202000.000000
Rwneg112_11 in112_11 sn112_11 78000.000000
Rwneg112_12 in112_12 sn112_12 78000.000000
Rwneg112_13 in112_13 sn112_13 202000.000000
Rwneg112_14 in112_14 sn112_14 202000.000000
Rwneg112_15 in112_15 sn112_15 202000.000000
Rwneg112_16 in112_16 sn112_16 202000.000000
Rwneg112_17 in112_17 sn112_17 78000.000000
Rwneg112_18 in112_18 sn112_18 202000.000000
Rwneg112_19 in112_19 sn112_19 78000.000000
Rwneg112_20 in112_20 sn112_20 202000.000000
Rwneg112_21 in112_21 sn112_21 202000.000000
Rwneg112_22 in112_22 sn112_22 78000.000000
Rwneg112_23 in112_23 sn112_23 202000.000000
Rwneg112_24 in112_24 sn112_24 78000.000000
Rwneg112_25 in112_25 sn112_25 202000.000000
Rwneg112_26 in112_26 sn112_26 202000.000000
Rwneg112_27 in112_27 sn112_27 78000.000000
Rwneg112_28 in112_28 sn112_28 202000.000000
Rwneg112_29 in112_29 sn112_29 202000.000000
Rwneg112_30 in112_30 sn112_30 202000.000000
Rwneg112_31 in112_31 sn112_31 78000.000000
Rwneg112_32 in112_32 sn112_32 78000.000000
Rwneg112_33 in112_33 sn112_33 202000.000000
Rwneg112_34 in112_34 sn112_34 202000.000000
Rwneg112_35 in112_35 sn112_35 78000.000000
Rwneg112_36 in112_36 sn112_36 202000.000000
Rwneg112_37 in112_37 sn112_37 202000.000000
Rwneg112_38 in112_38 sn112_38 78000.000000
Rwneg112_39 in112_39 sn112_39 202000.000000
Rwneg112_40 in112_40 sn112_40 78000.000000
Rwneg112_41 in112_41 sn112_41 202000.000000
Rwneg112_42 in112_42 sn112_42 202000.000000
Rwneg112_43 in112_43 sn112_43 202000.000000
Rwneg112_44 in112_44 sn112_44 202000.000000
Rwneg112_45 in112_45 sn112_45 202000.000000
Rwneg112_46 in112_46 sn112_46 78000.000000
Rwneg112_47 in112_47 sn112_47 202000.000000
Rwneg112_48 in112_48 sn112_48 78000.000000
Rwneg112_49 in112_49 sn112_49 78000.000000
Rwneg112_50 in112_50 sn112_50 202000.000000
Rwneg112_51 in112_51 sn112_51 202000.000000
Rwneg112_52 in112_52 sn112_52 202000.000000
Rwneg112_53 in112_53 sn112_53 78000.000000
Rwneg112_54 in112_54 sn112_54 202000.000000
Rwneg112_55 in112_55 sn112_55 202000.000000
Rwneg112_56 in112_56 sn112_56 202000.000000
Rwneg112_57 in112_57 sn112_57 78000.000000
Rwneg112_58 in112_58 sn112_58 202000.000000
Rwneg112_59 in112_59 sn112_59 78000.000000
Rwneg112_60 in112_60 sn112_60 202000.000000
Rwneg112_61 in112_61 sn112_61 78000.000000
Rwneg112_62 in112_62 sn112_62 202000.000000
Rwneg112_63 in112_63 sn112_63 78000.000000
Rwneg112_64 in112_64 sn112_64 78000.000000
Rwneg112_65 in112_65 sn112_65 202000.000000
Rwneg112_66 in112_66 sn112_66 202000.000000
Rwneg112_67 in112_67 sn112_67 78000.000000
Rwneg112_68 in112_68 sn112_68 202000.000000
Rwneg112_69 in112_69 sn112_69 202000.000000
Rwneg112_70 in112_70 sn112_70 202000.000000
Rwneg112_71 in112_71 sn112_71 202000.000000
Rwneg112_72 in112_72 sn112_72 78000.000000
Rwneg112_73 in112_73 sn112_73 78000.000000
Rwneg112_74 in112_74 sn112_74 78000.000000
Rwneg112_75 in112_75 sn112_75 78000.000000
Rwneg112_76 in112_76 sn112_76 78000.000000
Rwneg112_77 in112_77 sn112_77 202000.000000
Rwneg112_78 in112_78 sn112_78 202000.000000
Rwneg112_79 in112_79 sn112_79 202000.000000
Rwneg112_80 in112_80 sn112_80 202000.000000
Rwneg112_81 in112_81 sn112_81 202000.000000
Rwneg112_82 in112_82 sn112_82 78000.000000
Rwneg112_83 in112_83 sn112_83 202000.000000
Rwneg112_84 in112_84 sn112_84 202000.000000
Rwneg113_1 in113_1 sn113_1 202000.000000
Rwneg113_2 in113_2 sn113_2 78000.000000
Rwneg113_3 in113_3 sn113_3 202000.000000
Rwneg113_4 in113_4 sn113_4 202000.000000
Rwneg113_5 in113_5 sn113_5 202000.000000
Rwneg113_6 in113_6 sn113_6 202000.000000
Rwneg113_7 in113_7 sn113_7 78000.000000
Rwneg113_8 in113_8 sn113_8 202000.000000
Rwneg113_9 in113_9 sn113_9 78000.000000
Rwneg113_10 in113_10 sn113_10 78000.000000
Rwneg113_11 in113_11 sn113_11 202000.000000
Rwneg113_12 in113_12 sn113_12 202000.000000
Rwneg113_13 in113_13 sn113_13 202000.000000
Rwneg113_14 in113_14 sn113_14 202000.000000
Rwneg113_15 in113_15 sn113_15 78000.000000
Rwneg113_16 in113_16 sn113_16 202000.000000
Rwneg113_17 in113_17 sn113_17 202000.000000
Rwneg113_18 in113_18 sn113_18 202000.000000
Rwneg113_19 in113_19 sn113_19 78000.000000
Rwneg113_20 in113_20 sn113_20 202000.000000
Rwneg113_21 in113_21 sn113_21 78000.000000
Rwneg113_22 in113_22 sn113_22 202000.000000
Rwneg113_23 in113_23 sn113_23 202000.000000
Rwneg113_24 in113_24 sn113_24 202000.000000
Rwneg113_25 in113_25 sn113_25 78000.000000
Rwneg113_26 in113_26 sn113_26 78000.000000
Rwneg113_27 in113_27 sn113_27 202000.000000
Rwneg113_28 in113_28 sn113_28 202000.000000
Rwneg113_29 in113_29 sn113_29 78000.000000
Rwneg113_30 in113_30 sn113_30 202000.000000
Rwneg113_31 in113_31 sn113_31 202000.000000
Rwneg113_32 in113_32 sn113_32 78000.000000
Rwneg113_33 in113_33 sn113_33 78000.000000
Rwneg113_34 in113_34 sn113_34 202000.000000
Rwneg113_35 in113_35 sn113_35 202000.000000
Rwneg113_36 in113_36 sn113_36 78000.000000
Rwneg113_37 in113_37 sn113_37 78000.000000
Rwneg113_38 in113_38 sn113_38 78000.000000
Rwneg113_39 in113_39 sn113_39 78000.000000
Rwneg113_40 in113_40 sn113_40 202000.000000
Rwneg113_41 in113_41 sn113_41 202000.000000
Rwneg113_42 in113_42 sn113_42 78000.000000
Rwneg113_43 in113_43 sn113_43 202000.000000
Rwneg113_44 in113_44 sn113_44 202000.000000
Rwneg113_45 in113_45 sn113_45 202000.000000
Rwneg113_46 in113_46 sn113_46 202000.000000
Rwneg113_47 in113_47 sn113_47 78000.000000
Rwneg113_48 in113_48 sn113_48 202000.000000
Rwneg113_49 in113_49 sn113_49 78000.000000
Rwneg113_50 in113_50 sn113_50 78000.000000
Rwneg113_51 in113_51 sn113_51 78000.000000
Rwneg113_52 in113_52 sn113_52 78000.000000
Rwneg113_53 in113_53 sn113_53 78000.000000
Rwneg113_54 in113_54 sn113_54 202000.000000
Rwneg113_55 in113_55 sn113_55 78000.000000
Rwneg113_56 in113_56 sn113_56 202000.000000
Rwneg113_57 in113_57 sn113_57 202000.000000
Rwneg113_58 in113_58 sn113_58 202000.000000
Rwneg113_59 in113_59 sn113_59 202000.000000
Rwneg113_60 in113_60 sn113_60 78000.000000
Rwneg113_61 in113_61 sn113_61 78000.000000
Rwneg113_62 in113_62 sn113_62 202000.000000
Rwneg113_63 in113_63 sn113_63 78000.000000
Rwneg113_64 in113_64 sn113_64 202000.000000
Rwneg113_65 in113_65 sn113_65 202000.000000
Rwneg113_66 in113_66 sn113_66 78000.000000
Rwneg113_67 in113_67 sn113_67 78000.000000
Rwneg113_68 in113_68 sn113_68 202000.000000
Rwneg113_69 in113_69 sn113_69 202000.000000
Rwneg113_70 in113_70 sn113_70 202000.000000
Rwneg113_71 in113_71 sn113_71 202000.000000
Rwneg113_72 in113_72 sn113_72 202000.000000
Rwneg113_73 in113_73 sn113_73 202000.000000
Rwneg113_74 in113_74 sn113_74 78000.000000
Rwneg113_75 in113_75 sn113_75 202000.000000
Rwneg113_76 in113_76 sn113_76 78000.000000
Rwneg113_77 in113_77 sn113_77 202000.000000
Rwneg113_78 in113_78 sn113_78 78000.000000
Rwneg113_79 in113_79 sn113_79 78000.000000
Rwneg113_80 in113_80 sn113_80 202000.000000
Rwneg113_81 in113_81 sn113_81 202000.000000
Rwneg113_82 in113_82 sn113_82 78000.000000
Rwneg113_83 in113_83 sn113_83 78000.000000
Rwneg113_84 in113_84 sn113_84 78000.000000
Rwneg114_1 in114_1 sn114_1 78000.000000
Rwneg114_2 in114_2 sn114_2 202000.000000
Rwneg114_3 in114_3 sn114_3 202000.000000
Rwneg114_4 in114_4 sn114_4 202000.000000
Rwneg114_5 in114_5 sn114_5 78000.000000
Rwneg114_6 in114_6 sn114_6 202000.000000
Rwneg114_7 in114_7 sn114_7 202000.000000
Rwneg114_8 in114_8 sn114_8 78000.000000
Rwneg114_9 in114_9 sn114_9 78000.000000
Rwneg114_10 in114_10 sn114_10 202000.000000
Rwneg114_11 in114_11 sn114_11 202000.000000
Rwneg114_12 in114_12 sn114_12 78000.000000
Rwneg114_13 in114_13 sn114_13 202000.000000
Rwneg114_14 in114_14 sn114_14 202000.000000
Rwneg114_15 in114_15 sn114_15 202000.000000
Rwneg114_16 in114_16 sn114_16 202000.000000
Rwneg114_17 in114_17 sn114_17 78000.000000
Rwneg114_18 in114_18 sn114_18 78000.000000
Rwneg114_19 in114_19 sn114_19 202000.000000
Rwneg114_20 in114_20 sn114_20 202000.000000
Rwneg114_21 in114_21 sn114_21 202000.000000
Rwneg114_22 in114_22 sn114_22 202000.000000
Rwneg114_23 in114_23 sn114_23 202000.000000
Rwneg114_24 in114_24 sn114_24 78000.000000
Rwneg114_25 in114_25 sn114_25 202000.000000
Rwneg114_26 in114_26 sn114_26 202000.000000
Rwneg114_27 in114_27 sn114_27 78000.000000
Rwneg114_28 in114_28 sn114_28 202000.000000
Rwneg114_29 in114_29 sn114_29 202000.000000
Rwneg114_30 in114_30 sn114_30 202000.000000
Rwneg114_31 in114_31 sn114_31 202000.000000
Rwneg114_32 in114_32 sn114_32 78000.000000
Rwneg114_33 in114_33 sn114_33 202000.000000
Rwneg114_34 in114_34 sn114_34 78000.000000
Rwneg114_35 in114_35 sn114_35 202000.000000
Rwneg114_36 in114_36 sn114_36 78000.000000
Rwneg114_37 in114_37 sn114_37 202000.000000
Rwneg114_38 in114_38 sn114_38 202000.000000
Rwneg114_39 in114_39 sn114_39 78000.000000
Rwneg114_40 in114_40 sn114_40 202000.000000
Rwneg114_41 in114_41 sn114_41 78000.000000
Rwneg114_42 in114_42 sn114_42 202000.000000
Rwneg114_43 in114_43 sn114_43 202000.000000
Rwneg114_44 in114_44 sn114_44 78000.000000
Rwneg114_45 in114_45 sn114_45 202000.000000
Rwneg114_46 in114_46 sn114_46 202000.000000
Rwneg114_47 in114_47 sn114_47 202000.000000
Rwneg114_48 in114_48 sn114_48 202000.000000
Rwneg114_49 in114_49 sn114_49 202000.000000
Rwneg114_50 in114_50 sn114_50 202000.000000
Rwneg114_51 in114_51 sn114_51 202000.000000
Rwneg114_52 in114_52 sn114_52 202000.000000
Rwneg114_53 in114_53 sn114_53 202000.000000
Rwneg114_54 in114_54 sn114_54 202000.000000
Rwneg114_55 in114_55 sn114_55 202000.000000
Rwneg114_56 in114_56 sn114_56 78000.000000
Rwneg114_57 in114_57 sn114_57 78000.000000
Rwneg114_58 in114_58 sn114_58 202000.000000
Rwneg114_59 in114_59 sn114_59 202000.000000
Rwneg114_60 in114_60 sn114_60 78000.000000
Rwneg114_61 in114_61 sn114_61 78000.000000
Rwneg114_62 in114_62 sn114_62 202000.000000
Rwneg114_63 in114_63 sn114_63 202000.000000
Rwneg114_64 in114_64 sn114_64 78000.000000
Rwneg114_65 in114_65 sn114_65 202000.000000
Rwneg114_66 in114_66 sn114_66 202000.000000
Rwneg114_67 in114_67 sn114_67 202000.000000
Rwneg114_68 in114_68 sn114_68 78000.000000
Rwneg114_69 in114_69 sn114_69 78000.000000
Rwneg114_70 in114_70 sn114_70 202000.000000
Rwneg114_71 in114_71 sn114_71 78000.000000
Rwneg114_72 in114_72 sn114_72 202000.000000
Rwneg114_73 in114_73 sn114_73 78000.000000
Rwneg114_74 in114_74 sn114_74 78000.000000
Rwneg114_75 in114_75 sn114_75 78000.000000
Rwneg114_76 in114_76 sn114_76 202000.000000
Rwneg114_77 in114_77 sn114_77 78000.000000
Rwneg114_78 in114_78 sn114_78 78000.000000
Rwneg114_79 in114_79 sn114_79 78000.000000
Rwneg114_80 in114_80 sn114_80 78000.000000
Rwneg114_81 in114_81 sn114_81 202000.000000
Rwneg114_82 in114_82 sn114_82 78000.000000
Rwneg114_83 in114_83 sn114_83 78000.000000
Rwneg114_84 in114_84 sn114_84 202000.000000
Rwneg115_1 in115_1 sn115_1 202000.000000
Rwneg115_2 in115_2 sn115_2 202000.000000
Rwneg115_3 in115_3 sn115_3 202000.000000
Rwneg115_4 in115_4 sn115_4 78000.000000
Rwneg115_5 in115_5 sn115_5 202000.000000
Rwneg115_6 in115_6 sn115_6 202000.000000
Rwneg115_7 in115_7 sn115_7 78000.000000
Rwneg115_8 in115_8 sn115_8 202000.000000
Rwneg115_9 in115_9 sn115_9 202000.000000
Rwneg115_10 in115_10 sn115_10 78000.000000
Rwneg115_11 in115_11 sn115_11 202000.000000
Rwneg115_12 in115_12 sn115_12 78000.000000
Rwneg115_13 in115_13 sn115_13 78000.000000
Rwneg115_14 in115_14 sn115_14 78000.000000
Rwneg115_15 in115_15 sn115_15 202000.000000
Rwneg115_16 in115_16 sn115_16 78000.000000
Rwneg115_17 in115_17 sn115_17 202000.000000
Rwneg115_18 in115_18 sn115_18 78000.000000
Rwneg115_19 in115_19 sn115_19 202000.000000
Rwneg115_20 in115_20 sn115_20 78000.000000
Rwneg115_21 in115_21 sn115_21 202000.000000
Rwneg115_22 in115_22 sn115_22 202000.000000
Rwneg115_23 in115_23 sn115_23 78000.000000
Rwneg115_24 in115_24 sn115_24 202000.000000
Rwneg115_25 in115_25 sn115_25 202000.000000
Rwneg115_26 in115_26 sn115_26 78000.000000
Rwneg115_27 in115_27 sn115_27 202000.000000
Rwneg115_28 in115_28 sn115_28 78000.000000
Rwneg115_29 in115_29 sn115_29 202000.000000
Rwneg115_30 in115_30 sn115_30 202000.000000
Rwneg115_31 in115_31 sn115_31 202000.000000
Rwneg115_32 in115_32 sn115_32 78000.000000
Rwneg115_33 in115_33 sn115_33 202000.000000
Rwneg115_34 in115_34 sn115_34 78000.000000
Rwneg115_35 in115_35 sn115_35 78000.000000
Rwneg115_36 in115_36 sn115_36 202000.000000
Rwneg115_37 in115_37 sn115_37 78000.000000
Rwneg115_38 in115_38 sn115_38 78000.000000
Rwneg115_39 in115_39 sn115_39 78000.000000
Rwneg115_40 in115_40 sn115_40 78000.000000
Rwneg115_41 in115_41 sn115_41 78000.000000
Rwneg115_42 in115_42 sn115_42 78000.000000
Rwneg115_43 in115_43 sn115_43 202000.000000
Rwneg115_44 in115_44 sn115_44 202000.000000
Rwneg115_45 in115_45 sn115_45 78000.000000
Rwneg115_46 in115_46 sn115_46 202000.000000
Rwneg115_47 in115_47 sn115_47 78000.000000
Rwneg115_48 in115_48 sn115_48 78000.000000
Rwneg115_49 in115_49 sn115_49 78000.000000
Rwneg115_50 in115_50 sn115_50 78000.000000
Rwneg115_51 in115_51 sn115_51 78000.000000
Rwneg115_52 in115_52 sn115_52 78000.000000
Rwneg115_53 in115_53 sn115_53 202000.000000
Rwneg115_54 in115_54 sn115_54 202000.000000
Rwneg115_55 in115_55 sn115_55 78000.000000
Rwneg115_56 in115_56 sn115_56 202000.000000
Rwneg115_57 in115_57 sn115_57 202000.000000
Rwneg115_58 in115_58 sn115_58 202000.000000
Rwneg115_59 in115_59 sn115_59 202000.000000
Rwneg115_60 in115_60 sn115_60 202000.000000
Rwneg115_61 in115_61 sn115_61 202000.000000
Rwneg115_62 in115_62 sn115_62 78000.000000
Rwneg115_63 in115_63 sn115_63 78000.000000
Rwneg115_64 in115_64 sn115_64 202000.000000
Rwneg115_65 in115_65 sn115_65 202000.000000
Rwneg115_66 in115_66 sn115_66 202000.000000
Rwneg115_67 in115_67 sn115_67 202000.000000
Rwneg115_68 in115_68 sn115_68 78000.000000
Rwneg115_69 in115_69 sn115_69 78000.000000
Rwneg115_70 in115_70 sn115_70 78000.000000
Rwneg115_71 in115_71 sn115_71 78000.000000
Rwneg115_72 in115_72 sn115_72 78000.000000
Rwneg115_73 in115_73 sn115_73 202000.000000
Rwneg115_74 in115_74 sn115_74 202000.000000
Rwneg115_75 in115_75 sn115_75 78000.000000
Rwneg115_76 in115_76 sn115_76 202000.000000
Rwneg115_77 in115_77 sn115_77 78000.000000
Rwneg115_78 in115_78 sn115_78 202000.000000
Rwneg115_79 in115_79 sn115_79 78000.000000
Rwneg115_80 in115_80 sn115_80 78000.000000
Rwneg115_81 in115_81 sn115_81 78000.000000
Rwneg115_82 in115_82 sn115_82 202000.000000
Rwneg115_83 in115_83 sn115_83 202000.000000
Rwneg115_84 in115_84 sn115_84 78000.000000
Rwneg116_1 in116_1 sn116_1 202000.000000
Rwneg116_2 in116_2 sn116_2 78000.000000
Rwneg116_3 in116_3 sn116_3 78000.000000
Rwneg116_4 in116_4 sn116_4 202000.000000
Rwneg116_5 in116_5 sn116_5 202000.000000
Rwneg116_6 in116_6 sn116_6 78000.000000
Rwneg116_7 in116_7 sn116_7 78000.000000
Rwneg116_8 in116_8 sn116_8 78000.000000
Rwneg116_9 in116_9 sn116_9 202000.000000
Rwneg116_10 in116_10 sn116_10 78000.000000
Rwneg116_11 in116_11 sn116_11 202000.000000
Rwneg116_12 in116_12 sn116_12 202000.000000
Rwneg116_13 in116_13 sn116_13 78000.000000
Rwneg116_14 in116_14 sn116_14 202000.000000
Rwneg116_15 in116_15 sn116_15 202000.000000
Rwneg116_16 in116_16 sn116_16 78000.000000
Rwneg116_17 in116_17 sn116_17 78000.000000
Rwneg116_18 in116_18 sn116_18 202000.000000
Rwneg116_19 in116_19 sn116_19 78000.000000
Rwneg116_20 in116_20 sn116_20 78000.000000
Rwneg116_21 in116_21 sn116_21 78000.000000
Rwneg116_22 in116_22 sn116_22 78000.000000
Rwneg116_23 in116_23 sn116_23 202000.000000
Rwneg116_24 in116_24 sn116_24 78000.000000
Rwneg116_25 in116_25 sn116_25 78000.000000
Rwneg116_26 in116_26 sn116_26 78000.000000
Rwneg116_27 in116_27 sn116_27 78000.000000
Rwneg116_28 in116_28 sn116_28 202000.000000
Rwneg116_29 in116_29 sn116_29 202000.000000
Rwneg116_30 in116_30 sn116_30 78000.000000
Rwneg116_31 in116_31 sn116_31 202000.000000
Rwneg116_32 in116_32 sn116_32 202000.000000
Rwneg116_33 in116_33 sn116_33 78000.000000
Rwneg116_34 in116_34 sn116_34 202000.000000
Rwneg116_35 in116_35 sn116_35 202000.000000
Rwneg116_36 in116_36 sn116_36 202000.000000
Rwneg116_37 in116_37 sn116_37 202000.000000
Rwneg116_38 in116_38 sn116_38 78000.000000
Rwneg116_39 in116_39 sn116_39 202000.000000
Rwneg116_40 in116_40 sn116_40 202000.000000
Rwneg116_41 in116_41 sn116_41 78000.000000
Rwneg116_42 in116_42 sn116_42 78000.000000
Rwneg116_43 in116_43 sn116_43 202000.000000
Rwneg116_44 in116_44 sn116_44 78000.000000
Rwneg116_45 in116_45 sn116_45 78000.000000
Rwneg116_46 in116_46 sn116_46 202000.000000
Rwneg116_47 in116_47 sn116_47 202000.000000
Rwneg116_48 in116_48 sn116_48 78000.000000
Rwneg116_49 in116_49 sn116_49 202000.000000
Rwneg116_50 in116_50 sn116_50 202000.000000
Rwneg116_51 in116_51 sn116_51 202000.000000
Rwneg116_52 in116_52 sn116_52 202000.000000
Rwneg116_53 in116_53 sn116_53 202000.000000
Rwneg116_54 in116_54 sn116_54 78000.000000
Rwneg116_55 in116_55 sn116_55 202000.000000
Rwneg116_56 in116_56 sn116_56 202000.000000
Rwneg116_57 in116_57 sn116_57 202000.000000
Rwneg116_58 in116_58 sn116_58 202000.000000
Rwneg116_59 in116_59 sn116_59 202000.000000
Rwneg116_60 in116_60 sn116_60 78000.000000
Rwneg116_61 in116_61 sn116_61 202000.000000
Rwneg116_62 in116_62 sn116_62 202000.000000
Rwneg116_63 in116_63 sn116_63 78000.000000
Rwneg116_64 in116_64 sn116_64 78000.000000
Rwneg116_65 in116_65 sn116_65 78000.000000
Rwneg116_66 in116_66 sn116_66 202000.000000
Rwneg116_67 in116_67 sn116_67 202000.000000
Rwneg116_68 in116_68 sn116_68 202000.000000
Rwneg116_69 in116_69 sn116_69 202000.000000
Rwneg116_70 in116_70 sn116_70 78000.000000
Rwneg116_71 in116_71 sn116_71 202000.000000
Rwneg116_72 in116_72 sn116_72 78000.000000
Rwneg116_73 in116_73 sn116_73 202000.000000
Rwneg116_74 in116_74 sn116_74 78000.000000
Rwneg116_75 in116_75 sn116_75 202000.000000
Rwneg116_76 in116_76 sn116_76 202000.000000
Rwneg116_77 in116_77 sn116_77 202000.000000
Rwneg116_78 in116_78 sn116_78 202000.000000
Rwneg116_79 in116_79 sn116_79 202000.000000
Rwneg116_80 in116_80 sn116_80 202000.000000
Rwneg116_81 in116_81 sn116_81 78000.000000
Rwneg116_82 in116_82 sn116_82 202000.000000
Rwneg116_83 in116_83 sn116_83 78000.000000
Rwneg116_84 in116_84 sn116_84 78000.000000
Rwneg117_1 in117_1 sn117_1 202000.000000
Rwneg117_2 in117_2 sn117_2 202000.000000
Rwneg117_3 in117_3 sn117_3 78000.000000
Rwneg117_4 in117_4 sn117_4 78000.000000
Rwneg117_5 in117_5 sn117_5 202000.000000
Rwneg117_6 in117_6 sn117_6 78000.000000
Rwneg117_7 in117_7 sn117_7 202000.000000
Rwneg117_8 in117_8 sn117_8 202000.000000
Rwneg117_9 in117_9 sn117_9 202000.000000
Rwneg117_10 in117_10 sn117_10 202000.000000
Rwneg117_11 in117_11 sn117_11 78000.000000
Rwneg117_12 in117_12 sn117_12 202000.000000
Rwneg117_13 in117_13 sn117_13 202000.000000
Rwneg117_14 in117_14 sn117_14 78000.000000
Rwneg117_15 in117_15 sn117_15 78000.000000
Rwneg117_16 in117_16 sn117_16 202000.000000
Rwneg117_17 in117_17 sn117_17 78000.000000
Rwneg117_18 in117_18 sn117_18 78000.000000
Rwneg117_19 in117_19 sn117_19 78000.000000
Rwneg117_20 in117_20 sn117_20 202000.000000
Rwneg117_21 in117_21 sn117_21 202000.000000
Rwneg117_22 in117_22 sn117_22 78000.000000
Rwneg117_23 in117_23 sn117_23 78000.000000
Rwneg117_24 in117_24 sn117_24 78000.000000
Rwneg117_25 in117_25 sn117_25 202000.000000
Rwneg117_26 in117_26 sn117_26 202000.000000
Rwneg117_27 in117_27 sn117_27 202000.000000
Rwneg117_28 in117_28 sn117_28 202000.000000
Rwneg117_29 in117_29 sn117_29 78000.000000
Rwneg117_30 in117_30 sn117_30 202000.000000
Rwneg117_31 in117_31 sn117_31 78000.000000
Rwneg117_32 in117_32 sn117_32 202000.000000
Rwneg117_33 in117_33 sn117_33 202000.000000
Rwneg117_34 in117_34 sn117_34 78000.000000
Rwneg117_35 in117_35 sn117_35 202000.000000
Rwneg117_36 in117_36 sn117_36 78000.000000
Rwneg117_37 in117_37 sn117_37 202000.000000
Rwneg117_38 in117_38 sn117_38 78000.000000
Rwneg117_39 in117_39 sn117_39 78000.000000
Rwneg117_40 in117_40 sn117_40 78000.000000
Rwneg117_41 in117_41 sn117_41 78000.000000
Rwneg117_42 in117_42 sn117_42 202000.000000
Rwneg117_43 in117_43 sn117_43 202000.000000
Rwneg117_44 in117_44 sn117_44 202000.000000
Rwneg117_45 in117_45 sn117_45 202000.000000
Rwneg117_46 in117_46 sn117_46 78000.000000
Rwneg117_47 in117_47 sn117_47 202000.000000
Rwneg117_48 in117_48 sn117_48 78000.000000
Rwneg117_49 in117_49 sn117_49 78000.000000
Rwneg117_50 in117_50 sn117_50 202000.000000
Rwneg117_51 in117_51 sn117_51 202000.000000
Rwneg117_52 in117_52 sn117_52 202000.000000
Rwneg117_53 in117_53 sn117_53 78000.000000
Rwneg117_54 in117_54 sn117_54 202000.000000
Rwneg117_55 in117_55 sn117_55 202000.000000
Rwneg117_56 in117_56 sn117_56 78000.000000
Rwneg117_57 in117_57 sn117_57 78000.000000
Rwneg117_58 in117_58 sn117_58 78000.000000
Rwneg117_59 in117_59 sn117_59 202000.000000
Rwneg117_60 in117_60 sn117_60 202000.000000
Rwneg117_61 in117_61 sn117_61 202000.000000
Rwneg117_62 in117_62 sn117_62 202000.000000
Rwneg117_63 in117_63 sn117_63 202000.000000
Rwneg117_64 in117_64 sn117_64 202000.000000
Rwneg117_65 in117_65 sn117_65 78000.000000
Rwneg117_66 in117_66 sn117_66 202000.000000
Rwneg117_67 in117_67 sn117_67 78000.000000
Rwneg117_68 in117_68 sn117_68 78000.000000
Rwneg117_69 in117_69 sn117_69 202000.000000
Rwneg117_70 in117_70 sn117_70 78000.000000
Rwneg117_71 in117_71 sn117_71 78000.000000
Rwneg117_72 in117_72 sn117_72 202000.000000
Rwneg117_73 in117_73 sn117_73 202000.000000
Rwneg117_74 in117_74 sn117_74 202000.000000
Rwneg117_75 in117_75 sn117_75 78000.000000
Rwneg117_76 in117_76 sn117_76 202000.000000
Rwneg117_77 in117_77 sn117_77 78000.000000
Rwneg117_78 in117_78 sn117_78 78000.000000
Rwneg117_79 in117_79 sn117_79 78000.000000
Rwneg117_80 in117_80 sn117_80 202000.000000
Rwneg117_81 in117_81 sn117_81 202000.000000
Rwneg117_82 in117_82 sn117_82 202000.000000
Rwneg117_83 in117_83 sn117_83 202000.000000
Rwneg117_84 in117_84 sn117_84 78000.000000
Rwneg118_1 in118_1 sn118_1 78000.000000
Rwneg118_2 in118_2 sn118_2 78000.000000
Rwneg118_3 in118_3 sn118_3 202000.000000
Rwneg118_4 in118_4 sn118_4 202000.000000
Rwneg118_5 in118_5 sn118_5 202000.000000
Rwneg118_6 in118_6 sn118_6 202000.000000
Rwneg118_7 in118_7 sn118_7 78000.000000
Rwneg118_8 in118_8 sn118_8 78000.000000
Rwneg118_9 in118_9 sn118_9 78000.000000
Rwneg118_10 in118_10 sn118_10 202000.000000
Rwneg118_11 in118_11 sn118_11 202000.000000
Rwneg118_12 in118_12 sn118_12 202000.000000
Rwneg118_13 in118_13 sn118_13 202000.000000
Rwneg118_14 in118_14 sn118_14 202000.000000
Rwneg118_15 in118_15 sn118_15 78000.000000
Rwneg118_16 in118_16 sn118_16 202000.000000
Rwneg118_17 in118_17 sn118_17 202000.000000
Rwneg118_18 in118_18 sn118_18 202000.000000
Rwneg118_19 in118_19 sn118_19 202000.000000
Rwneg118_20 in118_20 sn118_20 202000.000000
Rwneg118_21 in118_21 sn118_21 202000.000000
Rwneg118_22 in118_22 sn118_22 78000.000000
Rwneg118_23 in118_23 sn118_23 202000.000000
Rwneg118_24 in118_24 sn118_24 78000.000000
Rwneg118_25 in118_25 sn118_25 78000.000000
Rwneg118_26 in118_26 sn118_26 78000.000000
Rwneg118_27 in118_27 sn118_27 78000.000000
Rwneg118_28 in118_28 sn118_28 78000.000000
Rwneg118_29 in118_29 sn118_29 202000.000000
Rwneg118_30 in118_30 sn118_30 78000.000000
Rwneg118_31 in118_31 sn118_31 202000.000000
Rwneg118_32 in118_32 sn118_32 202000.000000
Rwneg118_33 in118_33 sn118_33 202000.000000
Rwneg118_34 in118_34 sn118_34 202000.000000
Rwneg118_35 in118_35 sn118_35 78000.000000
Rwneg118_36 in118_36 sn118_36 78000.000000
Rwneg118_37 in118_37 sn118_37 202000.000000
Rwneg118_38 in118_38 sn118_38 202000.000000
Rwneg118_39 in118_39 sn118_39 78000.000000
Rwneg118_40 in118_40 sn118_40 202000.000000
Rwneg118_41 in118_41 sn118_41 78000.000000
Rwneg118_42 in118_42 sn118_42 78000.000000
Rwneg118_43 in118_43 sn118_43 202000.000000
Rwneg118_44 in118_44 sn118_44 78000.000000
Rwneg118_45 in118_45 sn118_45 202000.000000
Rwneg118_46 in118_46 sn118_46 202000.000000
Rwneg118_47 in118_47 sn118_47 78000.000000
Rwneg118_48 in118_48 sn118_48 202000.000000
Rwneg118_49 in118_49 sn118_49 78000.000000
Rwneg118_50 in118_50 sn118_50 202000.000000
Rwneg118_51 in118_51 sn118_51 202000.000000
Rwneg118_52 in118_52 sn118_52 78000.000000
Rwneg118_53 in118_53 sn118_53 202000.000000
Rwneg118_54 in118_54 sn118_54 78000.000000
Rwneg118_55 in118_55 sn118_55 78000.000000
Rwneg118_56 in118_56 sn118_56 202000.000000
Rwneg118_57 in118_57 sn118_57 78000.000000
Rwneg118_58 in118_58 sn118_58 202000.000000
Rwneg118_59 in118_59 sn118_59 202000.000000
Rwneg118_60 in118_60 sn118_60 78000.000000
Rwneg118_61 in118_61 sn118_61 202000.000000
Rwneg118_62 in118_62 sn118_62 202000.000000
Rwneg118_63 in118_63 sn118_63 78000.000000
Rwneg118_64 in118_64 sn118_64 202000.000000
Rwneg118_65 in118_65 sn118_65 78000.000000
Rwneg118_66 in118_66 sn118_66 202000.000000
Rwneg118_67 in118_67 sn118_67 202000.000000
Rwneg118_68 in118_68 sn118_68 202000.000000
Rwneg118_69 in118_69 sn118_69 202000.000000
Rwneg118_70 in118_70 sn118_70 78000.000000
Rwneg118_71 in118_71 sn118_71 202000.000000
Rwneg118_72 in118_72 sn118_72 78000.000000
Rwneg118_73 in118_73 sn118_73 202000.000000
Rwneg118_74 in118_74 sn118_74 78000.000000
Rwneg118_75 in118_75 sn118_75 202000.000000
Rwneg118_76 in118_76 sn118_76 78000.000000
Rwneg118_77 in118_77 sn118_77 202000.000000
Rwneg118_78 in118_78 sn118_78 78000.000000
Rwneg118_79 in118_79 sn118_79 202000.000000
Rwneg118_80 in118_80 sn118_80 202000.000000
Rwneg118_81 in118_81 sn118_81 202000.000000
Rwneg118_82 in118_82 sn118_82 78000.000000
Rwneg118_83 in118_83 sn118_83 202000.000000
Rwneg118_84 in118_84 sn118_84 202000.000000
Rwneg119_1 in119_1 sn119_1 78000.000000
Rwneg119_2 in119_2 sn119_2 202000.000000
Rwneg119_3 in119_3 sn119_3 78000.000000
Rwneg119_4 in119_4 sn119_4 78000.000000
Rwneg119_5 in119_5 sn119_5 78000.000000
Rwneg119_6 in119_6 sn119_6 78000.000000
Rwneg119_7 in119_7 sn119_7 202000.000000
Rwneg119_8 in119_8 sn119_8 78000.000000
Rwneg119_9 in119_9 sn119_9 202000.000000
Rwneg119_10 in119_10 sn119_10 78000.000000
Rwneg119_11 in119_11 sn119_11 202000.000000
Rwneg119_12 in119_12 sn119_12 78000.000000
Rwneg119_13 in119_13 sn119_13 78000.000000
Rwneg119_14 in119_14 sn119_14 78000.000000
Rwneg119_15 in119_15 sn119_15 202000.000000
Rwneg119_16 in119_16 sn119_16 202000.000000
Rwneg119_17 in119_17 sn119_17 202000.000000
Rwneg119_18 in119_18 sn119_18 78000.000000
Rwneg119_19 in119_19 sn119_19 202000.000000
Rwneg119_20 in119_20 sn119_20 78000.000000
Rwneg119_21 in119_21 sn119_21 202000.000000
Rwneg119_22 in119_22 sn119_22 202000.000000
Rwneg119_23 in119_23 sn119_23 202000.000000
Rwneg119_24 in119_24 sn119_24 202000.000000
Rwneg119_25 in119_25 sn119_25 202000.000000
Rwneg119_26 in119_26 sn119_26 78000.000000
Rwneg119_27 in119_27 sn119_27 78000.000000
Rwneg119_28 in119_28 sn119_28 78000.000000
Rwneg119_29 in119_29 sn119_29 202000.000000
Rwneg119_30 in119_30 sn119_30 202000.000000
Rwneg119_31 in119_31 sn119_31 78000.000000
Rwneg119_32 in119_32 sn119_32 202000.000000
Rwneg119_33 in119_33 sn119_33 78000.000000
Rwneg119_34 in119_34 sn119_34 202000.000000
Rwneg119_35 in119_35 sn119_35 78000.000000
Rwneg119_36 in119_36 sn119_36 202000.000000
Rwneg119_37 in119_37 sn119_37 202000.000000
Rwneg119_38 in119_38 sn119_38 202000.000000
Rwneg119_39 in119_39 sn119_39 78000.000000
Rwneg119_40 in119_40 sn119_40 202000.000000
Rwneg119_41 in119_41 sn119_41 202000.000000
Rwneg119_42 in119_42 sn119_42 78000.000000
Rwneg119_43 in119_43 sn119_43 202000.000000
Rwneg119_44 in119_44 sn119_44 202000.000000
Rwneg119_45 in119_45 sn119_45 202000.000000
Rwneg119_46 in119_46 sn119_46 78000.000000
Rwneg119_47 in119_47 sn119_47 78000.000000
Rwneg119_48 in119_48 sn119_48 202000.000000
Rwneg119_49 in119_49 sn119_49 202000.000000
Rwneg119_50 in119_50 sn119_50 202000.000000
Rwneg119_51 in119_51 sn119_51 78000.000000
Rwneg119_52 in119_52 sn119_52 202000.000000
Rwneg119_53 in119_53 sn119_53 78000.000000
Rwneg119_54 in119_54 sn119_54 78000.000000
Rwneg119_55 in119_55 sn119_55 78000.000000
Rwneg119_56 in119_56 sn119_56 202000.000000
Rwneg119_57 in119_57 sn119_57 202000.000000
Rwneg119_58 in119_58 sn119_58 202000.000000
Rwneg119_59 in119_59 sn119_59 78000.000000
Rwneg119_60 in119_60 sn119_60 202000.000000
Rwneg119_61 in119_61 sn119_61 202000.000000
Rwneg119_62 in119_62 sn119_62 78000.000000
Rwneg119_63 in119_63 sn119_63 78000.000000
Rwneg119_64 in119_64 sn119_64 202000.000000
Rwneg119_65 in119_65 sn119_65 202000.000000
Rwneg119_66 in119_66 sn119_66 78000.000000
Rwneg119_67 in119_67 sn119_67 78000.000000
Rwneg119_68 in119_68 sn119_68 202000.000000
Rwneg119_69 in119_69 sn119_69 78000.000000
Rwneg119_70 in119_70 sn119_70 78000.000000
Rwneg119_71 in119_71 sn119_71 78000.000000
Rwneg119_72 in119_72 sn119_72 202000.000000
Rwneg119_73 in119_73 sn119_73 202000.000000
Rwneg119_74 in119_74 sn119_74 202000.000000
Rwneg119_75 in119_75 sn119_75 78000.000000
Rwneg119_76 in119_76 sn119_76 78000.000000
Rwneg119_77 in119_77 sn119_77 202000.000000
Rwneg119_78 in119_78 sn119_78 202000.000000
Rwneg119_79 in119_79 sn119_79 202000.000000
Rwneg119_80 in119_80 sn119_80 78000.000000
Rwneg119_81 in119_81 sn119_81 78000.000000
Rwneg119_82 in119_82 sn119_82 202000.000000
Rwneg119_83 in119_83 sn119_83 202000.000000
Rwneg119_84 in119_84 sn119_84 78000.000000
Rwneg120_1 in120_1 sn120_1 202000.000000
Rwneg120_2 in120_2 sn120_2 78000.000000
Rwneg120_3 in120_3 sn120_3 202000.000000
Rwneg120_4 in120_4 sn120_4 202000.000000
Rwneg120_5 in120_5 sn120_5 202000.000000
Rwneg120_6 in120_6 sn120_6 78000.000000
Rwneg120_7 in120_7 sn120_7 78000.000000
Rwneg120_8 in120_8 sn120_8 78000.000000
Rwneg120_9 in120_9 sn120_9 78000.000000
Rwneg120_10 in120_10 sn120_10 78000.000000
Rwneg120_11 in120_11 sn120_11 202000.000000
Rwneg120_12 in120_12 sn120_12 78000.000000
Rwneg120_13 in120_13 sn120_13 202000.000000
Rwneg120_14 in120_14 sn120_14 202000.000000
Rwneg120_15 in120_15 sn120_15 78000.000000
Rwneg120_16 in120_16 sn120_16 202000.000000
Rwneg120_17 in120_17 sn120_17 202000.000000
Rwneg120_18 in120_18 sn120_18 78000.000000
Rwneg120_19 in120_19 sn120_19 202000.000000
Rwneg120_20 in120_20 sn120_20 78000.000000
Rwneg120_21 in120_21 sn120_21 202000.000000
Rwneg120_22 in120_22 sn120_22 202000.000000
Rwneg120_23 in120_23 sn120_23 78000.000000
Rwneg120_24 in120_24 sn120_24 78000.000000
Rwneg120_25 in120_25 sn120_25 202000.000000
Rwneg120_26 in120_26 sn120_26 78000.000000
Rwneg120_27 in120_27 sn120_27 202000.000000
Rwneg120_28 in120_28 sn120_28 202000.000000
Rwneg120_29 in120_29 sn120_29 78000.000000
Rwneg120_30 in120_30 sn120_30 202000.000000
Rwneg120_31 in120_31 sn120_31 202000.000000
Rwneg120_32 in120_32 sn120_32 202000.000000
Rwneg120_33 in120_33 sn120_33 202000.000000
Rwneg120_34 in120_34 sn120_34 78000.000000
Rwneg120_35 in120_35 sn120_35 202000.000000
Rwneg120_36 in120_36 sn120_36 78000.000000
Rwneg120_37 in120_37 sn120_37 78000.000000
Rwneg120_38 in120_38 sn120_38 202000.000000
Rwneg120_39 in120_39 sn120_39 78000.000000
Rwneg120_40 in120_40 sn120_40 78000.000000
Rwneg120_41 in120_41 sn120_41 78000.000000
Rwneg120_42 in120_42 sn120_42 78000.000000
Rwneg120_43 in120_43 sn120_43 202000.000000
Rwneg120_44 in120_44 sn120_44 202000.000000
Rwneg120_45 in120_45 sn120_45 78000.000000
Rwneg120_46 in120_46 sn120_46 78000.000000
Rwneg120_47 in120_47 sn120_47 78000.000000
Rwneg120_48 in120_48 sn120_48 78000.000000
Rwneg120_49 in120_49 sn120_49 78000.000000
Rwneg120_50 in120_50 sn120_50 78000.000000
Rwneg120_51 in120_51 sn120_51 78000.000000
Rwneg120_52 in120_52 sn120_52 78000.000000
Rwneg120_53 in120_53 sn120_53 78000.000000
Rwneg120_54 in120_54 sn120_54 202000.000000
Rwneg120_55 in120_55 sn120_55 78000.000000
Rwneg120_56 in120_56 sn120_56 202000.000000
Rwneg120_57 in120_57 sn120_57 202000.000000
Rwneg120_58 in120_58 sn120_58 202000.000000
Rwneg120_59 in120_59 sn120_59 202000.000000
Rwneg120_60 in120_60 sn120_60 78000.000000
Rwneg120_61 in120_61 sn120_61 202000.000000
Rwneg120_62 in120_62 sn120_62 78000.000000
Rwneg120_63 in120_63 sn120_63 78000.000000
Rwneg120_64 in120_64 sn120_64 78000.000000
Rwneg120_65 in120_65 sn120_65 202000.000000
Rwneg120_66 in120_66 sn120_66 78000.000000
Rwneg120_67 in120_67 sn120_67 78000.000000
Rwneg120_68 in120_68 sn120_68 78000.000000
Rwneg120_69 in120_69 sn120_69 202000.000000
Rwneg120_70 in120_70 sn120_70 202000.000000
Rwneg120_71 in120_71 sn120_71 78000.000000
Rwneg120_72 in120_72 sn120_72 202000.000000
Rwneg120_73 in120_73 sn120_73 202000.000000
Rwneg120_74 in120_74 sn120_74 202000.000000
Rwneg120_75 in120_75 sn120_75 78000.000000
Rwneg120_76 in120_76 sn120_76 78000.000000
Rwneg120_77 in120_77 sn120_77 78000.000000
Rwneg120_78 in120_78 sn120_78 202000.000000
Rwneg120_79 in120_79 sn120_79 78000.000000
Rwneg120_80 in120_80 sn120_80 202000.000000
Rwneg120_81 in120_81 sn120_81 78000.000000
Rwneg120_82 in120_82 sn120_82 78000.000000
Rwneg120_83 in120_83 sn120_83 202000.000000
Rwneg120_84 in120_84 sn120_84 78000.000000


**********Positive Biases**********

Rbpos1 vd1 sp121_1 78000.000000
Rbpos2 vd2 sp121_2 78000.000000
Rbpos3 vd3 sp121_3 78000.000000
Rbpos4 vd4 sp121_4 78000.000000
Rbpos5 vd5 sp121_5 78000.000000
Rbpos6 vd6 sp121_6 202000.000000
Rbpos7 vd7 sp121_7 78000.000000
Rbpos8 vd8 sp121_8 78000.000000
Rbpos9 vd9 sp121_9 78000.000000
Rbpos10 vd10 sp121_10 78000.000000
Rbpos11 vd11 sp121_11 78000.000000
Rbpos12 vd12 sp121_12 78000.000000
Rbpos13 vd13 sp121_13 202000.000000
Rbpos14 vd14 sp121_14 78000.000000
Rbpos15 vd15 sp121_15 202000.000000
Rbpos16 vd16 sp121_16 202000.000000
Rbpos17 vd17 sp121_17 202000.000000
Rbpos18 vd18 sp121_18 78000.000000
Rbpos19 vd19 sp121_19 78000.000000
Rbpos20 vd20 sp121_20 78000.000000
Rbpos21 vd21 sp121_21 78000.000000
Rbpos22 vd22 sp121_22 78000.000000
Rbpos23 vd23 sp121_23 202000.000000
Rbpos24 vd24 sp121_24 202000.000000
Rbpos25 vd25 sp121_25 202000.000000
Rbpos26 vd26 sp121_26 78000.000000
Rbpos27 vd27 sp121_27 202000.000000
Rbpos28 vd28 sp121_28 202000.000000
Rbpos29 vd29 sp121_29 78000.000000
Rbpos30 vd30 sp121_30 78000.000000
Rbpos31 vd31 sp121_31 202000.000000
Rbpos32 vd32 sp121_32 78000.000000
Rbpos33 vd33 sp121_33 78000.000000
Rbpos34 vd34 sp121_34 78000.000000
Rbpos35 vd35 sp121_35 78000.000000
Rbpos36 vd36 sp121_36 78000.000000
Rbpos37 vd37 sp121_37 78000.000000
Rbpos38 vd38 sp121_38 78000.000000
Rbpos39 vd39 sp121_39 78000.000000
Rbpos40 vd40 sp121_40 78000.000000
Rbpos41 vd41 sp121_41 202000.000000
Rbpos42 vd42 sp121_42 202000.000000
Rbpos43 vd43 sp121_43 78000.000000
Rbpos44 vd44 sp121_44 78000.000000
Rbpos45 vd45 sp121_45 78000.000000
Rbpos46 vd46 sp121_46 78000.000000
Rbpos47 vd47 sp121_47 78000.000000
Rbpos48 vd48 sp121_48 202000.000000
Rbpos49 vd49 sp121_49 78000.000000
Rbpos50 vd50 sp121_50 78000.000000
Rbpos51 vd51 sp121_51 202000.000000
Rbpos52 vd52 sp121_52 202000.000000
Rbpos53 vd53 sp121_53 202000.000000
Rbpos54 vd54 sp121_54 202000.000000
Rbpos55 vd55 sp121_55 78000.000000
Rbpos56 vd56 sp121_56 78000.000000
Rbpos57 vd57 sp121_57 78000.000000
Rbpos58 vd58 sp121_58 202000.000000
Rbpos59 vd59 sp121_59 78000.000000
Rbpos60 vd60 sp121_60 78000.000000
Rbpos61 vd61 sp121_61 202000.000000
Rbpos62 vd62 sp121_62 202000.000000
Rbpos63 vd63 sp121_63 78000.000000
Rbpos64 vd64 sp121_64 202000.000000
Rbpos65 vd65 sp121_65 202000.000000
Rbpos66 vd66 sp121_66 78000.000000
Rbpos67 vd67 sp121_67 78000.000000
Rbpos68 vd68 sp121_68 78000.000000
Rbpos69 vd69 sp121_69 78000.000000
Rbpos70 vd70 sp121_70 78000.000000
Rbpos71 vd71 sp121_71 78000.000000
Rbpos72 vd72 sp121_72 202000.000000
Rbpos73 vd73 sp121_73 202000.000000
Rbpos74 vd74 sp121_74 78000.000000
Rbpos75 vd75 sp121_75 78000.000000
Rbpos76 vd76 sp121_76 78000.000000
Rbpos77 vd77 sp121_77 78000.000000
Rbpos78 vd78 sp121_78 78000.000000
Rbpos79 vd79 sp121_79 78000.000000
Rbpos80 vd80 sp121_80 78000.000000
Rbpos81 vd81 sp121_81 202000.000000
Rbpos82 vd82 sp121_82 78000.000000
Rbpos83 vd83 sp121_83 202000.000000
Rbpos84 vd84 sp121_84 78000.000000


**********Negative Biases**********

Rbneg1 vd1 sn121_1 202000.000000
Rbneg2 vd2 sn121_2 202000.000000
Rbneg3 vd3 sn121_3 202000.000000
Rbneg4 vd4 sn121_4 202000.000000
Rbneg5 vd5 sn121_5 202000.000000
Rbneg6 vd6 sn121_6 78000.000000
Rbneg7 vd7 sn121_7 202000.000000
Rbneg8 vd8 sn121_8 202000.000000
Rbneg9 vd9 sn121_9 202000.000000
Rbneg10 vd10 sn121_10 202000.000000
Rbneg11 vd11 sn121_11 202000.000000
Rbneg12 vd12 sn121_12 202000.000000
Rbneg13 vd13 sn121_13 78000.000000
Rbneg14 vd14 sn121_14 202000.000000
Rbneg15 vd15 sn121_15 78000.000000
Rbneg16 vd16 sn121_16 78000.000000
Rbneg17 vd17 sn121_17 78000.000000
Rbneg18 vd18 sn121_18 202000.000000
Rbneg19 vd19 sn121_19 202000.000000
Rbneg20 vd20 sn121_20 202000.000000
Rbneg21 vd21 sn121_21 202000.000000
Rbneg22 vd22 sn121_22 202000.000000
Rbneg23 vd23 sn121_23 78000.000000
Rbneg24 vd24 sn121_24 78000.000000
Rbneg25 vd25 sn121_25 78000.000000
Rbneg26 vd26 sn121_26 202000.000000
Rbneg27 vd27 sn121_27 78000.000000
Rbneg28 vd28 sn121_28 78000.000000
Rbneg29 vd29 sn121_29 202000.000000
Rbneg30 vd30 sn121_30 202000.000000
Rbneg31 vd31 sn121_31 78000.000000
Rbneg32 vd32 sn121_32 202000.000000
Rbneg33 vd33 sn121_33 202000.000000
Rbneg34 vd34 sn121_34 202000.000000
Rbneg35 vd35 sn121_35 202000.000000
Rbneg36 vd36 sn121_36 202000.000000
Rbneg37 vd37 sn121_37 202000.000000
Rbneg38 vd38 sn121_38 202000.000000
Rbneg39 vd39 sn121_39 202000.000000
Rbneg40 vd40 sn121_40 202000.000000
Rbneg41 vd41 sn121_41 78000.000000
Rbneg42 vd42 sn121_42 78000.000000
Rbneg43 vd43 sn121_43 202000.000000
Rbneg44 vd44 sn121_44 202000.000000
Rbneg45 vd45 sn121_45 202000.000000
Rbneg46 vd46 sn121_46 202000.000000
Rbneg47 vd47 sn121_47 202000.000000
Rbneg48 vd48 sn121_48 78000.000000
Rbneg49 vd49 sn121_49 202000.000000
Rbneg50 vd50 sn121_50 202000.000000
Rbneg51 vd51 sn121_51 78000.000000
Rbneg52 vd52 sn121_52 78000.000000
Rbneg53 vd53 sn121_53 78000.000000
Rbneg54 vd54 sn121_54 78000.000000
Rbneg55 vd55 sn121_55 202000.000000
Rbneg56 vd56 sn121_56 202000.000000
Rbneg57 vd57 sn121_57 202000.000000
Rbneg58 vd58 sn121_58 78000.000000
Rbneg59 vd59 sn121_59 202000.000000
Rbneg60 vd60 sn121_60 202000.000000
Rbneg61 vd61 sn121_61 78000.000000
Rbneg62 vd62 sn121_62 78000.000000
Rbneg63 vd63 sn121_63 202000.000000
Rbneg64 vd64 sn121_64 78000.000000
Rbneg65 vd65 sn121_65 78000.000000
Rbneg66 vd66 sn121_66 202000.000000
Rbneg67 vd67 sn121_67 202000.000000
Rbneg68 vd68 sn121_68 202000.000000
Rbneg69 vd69 sn121_69 202000.000000
Rbneg70 vd70 sn121_70 202000.000000
Rbneg71 vd71 sn121_71 202000.000000
Rbneg72 vd72 sn121_72 78000.000000
Rbneg73 vd73 sn121_73 78000.000000
Rbneg74 vd74 sn121_74 202000.000000
Rbneg75 vd75 sn121_75 202000.000000
Rbneg76 vd76 sn121_76 202000.000000
Rbneg77 vd77 sn121_77 202000.000000
Rbneg78 vd78 sn121_78 202000.000000
Rbneg79 vd79 sn121_79 202000.000000
Rbneg80 vd80 sn121_80 202000.000000
Rbneg81 vd81 sn121_81 78000.000000
Rbneg82 vd82 sn121_82 202000.000000
Rbneg83 vd83 sn121_83 78000.000000
Rbneg84 vd84 sn121_84 202000.000000


**********Parasitic Resistances for Vertical Lines**********

Rin1_1 in1 in1_1 9.241569
Rin1_2 in1_1 in1_2 9.241569
Rin1_3 in1_2 in1_3 9.241569
Rin1_4 in1_3 in1_4 9.241569
Rin1_5 in1_4 in1_5 9.241569
Rin1_6 in1_5 in1_6 9.241569
Rin1_7 in1_6 in1_7 9.241569
Rin1_8 in1_7 in1_8 9.241569
Rin1_9 in1_8 in1_9 9.241569
Rin1_10 in1_9 in1_10 9.241569
Rin1_11 in1_10 in1_11 9.241569
Rin1_12 in1_11 in1_12 9.241569
Rin1_13 in1_12 in1_13 9.241569
Rin1_14 in1_13 in1_14 9.241569
Rin1_15 in1_14 in1_15 9.241569
Rin1_16 in1_15 in1_16 9.241569
Rin1_17 in1_16 in1_17 9.241569
Rin1_18 in1_17 in1_18 9.241569
Rin1_19 in1_18 in1_19 9.241569
Rin1_20 in1_19 in1_20 9.241569
Rin1_21 in1_20 in1_21 9.241569
Rin1_22 in1_21 in1_22 9.241569
Rin1_23 in1_22 in1_23 9.241569
Rin1_24 in1_23 in1_24 9.241569
Rin1_25 in1_24 in1_25 9.241569
Rin1_26 in1_25 in1_26 9.241569
Rin1_27 in1_26 in1_27 9.241569
Rin1_28 in1_27 in1_28 9.241569
Rin1_29 in1 in1_29 9.241569
Rin1_30 in1_29 in1_30 9.241569
Rin1_31 in1_30 in1_31 9.241569
Rin1_32 in1_31 in1_32 9.241569
Rin1_33 in1_32 in1_33 9.241569
Rin1_34 in1_33 in1_34 9.241569
Rin1_35 in1_34 in1_35 9.241569
Rin1_36 in1_35 in1_36 9.241569
Rin1_37 in1_36 in1_37 9.241569
Rin1_38 in1_37 in1_38 9.241569
Rin1_39 in1_38 in1_39 9.241569
Rin1_40 in1_39 in1_40 9.241569
Rin1_41 in1_40 in1_41 9.241569
Rin1_42 in1_41 in1_42 9.241569
Rin1_43 in1_42 in1_43 9.241569
Rin1_44 in1_43 in1_44 9.241569
Rin1_45 in1_44 in1_45 9.241569
Rin1_46 in1_45 in1_46 9.241569
Rin1_47 in1_46 in1_47 9.241569
Rin1_48 in1_47 in1_48 9.241569
Rin1_49 in1_48 in1_49 9.241569
Rin1_50 in1_49 in1_50 9.241569
Rin1_51 in1_50 in1_51 9.241569
Rin1_52 in1_51 in1_52 9.241569
Rin1_53 in1_52 in1_53 9.241569
Rin1_54 in1_53 in1_54 9.241569
Rin1_55 in1_54 in1_55 9.241569
Rin1_56 in1_55 in1_56 9.241569
Rin1_57 in1 in1_57 9.241569
Rin1_58 in1_57 in1_58 9.241569
Rin1_59 in1_58 in1_59 9.241569
Rin1_60 in1_59 in1_60 9.241569
Rin1_61 in1_60 in1_61 9.241569
Rin1_62 in1_61 in1_62 9.241569
Rin1_63 in1_62 in1_63 9.241569
Rin1_64 in1_63 in1_64 9.241569
Rin1_65 in1_64 in1_65 9.241569
Rin1_66 in1_65 in1_66 9.241569
Rin1_67 in1_66 in1_67 9.241569
Rin1_68 in1_67 in1_68 9.241569
Rin1_69 in1_68 in1_69 9.241569
Rin1_70 in1_69 in1_70 9.241569
Rin1_71 in1_70 in1_71 9.241569
Rin1_72 in1_71 in1_72 9.241569
Rin1_73 in1_72 in1_73 9.241569
Rin1_74 in1_73 in1_74 9.241569
Rin1_75 in1_74 in1_75 9.241569
Rin1_76 in1_75 in1_76 9.241569
Rin1_77 in1_76 in1_77 9.241569
Rin1_78 in1_77 in1_78 9.241569
Rin1_79 in1_78 in1_79 9.241569
Rin1_80 in1_79 in1_80 9.241569
Rin1_81 in1_80 in1_81 9.241569
Rin1_82 in1_81 in1_82 9.241569
Rin1_83 in1_82 in1_83 9.241569
Rin1_84 in1_83 in1_84 9.241569
Rin2_1 in2 in2_1 9.241569
Rin2_2 in2_1 in2_2 9.241569
Rin2_3 in2_2 in2_3 9.241569
Rin2_4 in2_3 in2_4 9.241569
Rin2_5 in2_4 in2_5 9.241569
Rin2_6 in2_5 in2_6 9.241569
Rin2_7 in2_6 in2_7 9.241569
Rin2_8 in2_7 in2_8 9.241569
Rin2_9 in2_8 in2_9 9.241569
Rin2_10 in2_9 in2_10 9.241569
Rin2_11 in2_10 in2_11 9.241569
Rin2_12 in2_11 in2_12 9.241569
Rin2_13 in2_12 in2_13 9.241569
Rin2_14 in2_13 in2_14 9.241569
Rin2_15 in2_14 in2_15 9.241569
Rin2_16 in2_15 in2_16 9.241569
Rin2_17 in2_16 in2_17 9.241569
Rin2_18 in2_17 in2_18 9.241569
Rin2_19 in2_18 in2_19 9.241569
Rin2_20 in2_19 in2_20 9.241569
Rin2_21 in2_20 in2_21 9.241569
Rin2_22 in2_21 in2_22 9.241569
Rin2_23 in2_22 in2_23 9.241569
Rin2_24 in2_23 in2_24 9.241569
Rin2_25 in2_24 in2_25 9.241569
Rin2_26 in2_25 in2_26 9.241569
Rin2_27 in2_26 in2_27 9.241569
Rin2_28 in2_27 in2_28 9.241569
Rin2_29 in2 in2_29 9.241569
Rin2_30 in2_29 in2_30 9.241569
Rin2_31 in2_30 in2_31 9.241569
Rin2_32 in2_31 in2_32 9.241569
Rin2_33 in2_32 in2_33 9.241569
Rin2_34 in2_33 in2_34 9.241569
Rin2_35 in2_34 in2_35 9.241569
Rin2_36 in2_35 in2_36 9.241569
Rin2_37 in2_36 in2_37 9.241569
Rin2_38 in2_37 in2_38 9.241569
Rin2_39 in2_38 in2_39 9.241569
Rin2_40 in2_39 in2_40 9.241569
Rin2_41 in2_40 in2_41 9.241569
Rin2_42 in2_41 in2_42 9.241569
Rin2_43 in2_42 in2_43 9.241569
Rin2_44 in2_43 in2_44 9.241569
Rin2_45 in2_44 in2_45 9.241569
Rin2_46 in2_45 in2_46 9.241569
Rin2_47 in2_46 in2_47 9.241569
Rin2_48 in2_47 in2_48 9.241569
Rin2_49 in2_48 in2_49 9.241569
Rin2_50 in2_49 in2_50 9.241569
Rin2_51 in2_50 in2_51 9.241569
Rin2_52 in2_51 in2_52 9.241569
Rin2_53 in2_52 in2_53 9.241569
Rin2_54 in2_53 in2_54 9.241569
Rin2_55 in2_54 in2_55 9.241569
Rin2_56 in2_55 in2_56 9.241569
Rin2_57 in2 in2_57 9.241569
Rin2_58 in2_57 in2_58 9.241569
Rin2_59 in2_58 in2_59 9.241569
Rin2_60 in2_59 in2_60 9.241569
Rin2_61 in2_60 in2_61 9.241569
Rin2_62 in2_61 in2_62 9.241569
Rin2_63 in2_62 in2_63 9.241569
Rin2_64 in2_63 in2_64 9.241569
Rin2_65 in2_64 in2_65 9.241569
Rin2_66 in2_65 in2_66 9.241569
Rin2_67 in2_66 in2_67 9.241569
Rin2_68 in2_67 in2_68 9.241569
Rin2_69 in2_68 in2_69 9.241569
Rin2_70 in2_69 in2_70 9.241569
Rin2_71 in2_70 in2_71 9.241569
Rin2_72 in2_71 in2_72 9.241569
Rin2_73 in2_72 in2_73 9.241569
Rin2_74 in2_73 in2_74 9.241569
Rin2_75 in2_74 in2_75 9.241569
Rin2_76 in2_75 in2_76 9.241569
Rin2_77 in2_76 in2_77 9.241569
Rin2_78 in2_77 in2_78 9.241569
Rin2_79 in2_78 in2_79 9.241569
Rin2_80 in2_79 in2_80 9.241569
Rin2_81 in2_80 in2_81 9.241569
Rin2_82 in2_81 in2_82 9.241569
Rin2_83 in2_82 in2_83 9.241569
Rin2_84 in2_83 in2_84 9.241569
Rin3_1 in3 in3_1 9.241569
Rin3_2 in3_1 in3_2 9.241569
Rin3_3 in3_2 in3_3 9.241569
Rin3_4 in3_3 in3_4 9.241569
Rin3_5 in3_4 in3_5 9.241569
Rin3_6 in3_5 in3_6 9.241569
Rin3_7 in3_6 in3_7 9.241569
Rin3_8 in3_7 in3_8 9.241569
Rin3_9 in3_8 in3_9 9.241569
Rin3_10 in3_9 in3_10 9.241569
Rin3_11 in3_10 in3_11 9.241569
Rin3_12 in3_11 in3_12 9.241569
Rin3_13 in3_12 in3_13 9.241569
Rin3_14 in3_13 in3_14 9.241569
Rin3_15 in3_14 in3_15 9.241569
Rin3_16 in3_15 in3_16 9.241569
Rin3_17 in3_16 in3_17 9.241569
Rin3_18 in3_17 in3_18 9.241569
Rin3_19 in3_18 in3_19 9.241569
Rin3_20 in3_19 in3_20 9.241569
Rin3_21 in3_20 in3_21 9.241569
Rin3_22 in3_21 in3_22 9.241569
Rin3_23 in3_22 in3_23 9.241569
Rin3_24 in3_23 in3_24 9.241569
Rin3_25 in3_24 in3_25 9.241569
Rin3_26 in3_25 in3_26 9.241569
Rin3_27 in3_26 in3_27 9.241569
Rin3_28 in3_27 in3_28 9.241569
Rin3_29 in3 in3_29 9.241569
Rin3_30 in3_29 in3_30 9.241569
Rin3_31 in3_30 in3_31 9.241569
Rin3_32 in3_31 in3_32 9.241569
Rin3_33 in3_32 in3_33 9.241569
Rin3_34 in3_33 in3_34 9.241569
Rin3_35 in3_34 in3_35 9.241569
Rin3_36 in3_35 in3_36 9.241569
Rin3_37 in3_36 in3_37 9.241569
Rin3_38 in3_37 in3_38 9.241569
Rin3_39 in3_38 in3_39 9.241569
Rin3_40 in3_39 in3_40 9.241569
Rin3_41 in3_40 in3_41 9.241569
Rin3_42 in3_41 in3_42 9.241569
Rin3_43 in3_42 in3_43 9.241569
Rin3_44 in3_43 in3_44 9.241569
Rin3_45 in3_44 in3_45 9.241569
Rin3_46 in3_45 in3_46 9.241569
Rin3_47 in3_46 in3_47 9.241569
Rin3_48 in3_47 in3_48 9.241569
Rin3_49 in3_48 in3_49 9.241569
Rin3_50 in3_49 in3_50 9.241569
Rin3_51 in3_50 in3_51 9.241569
Rin3_52 in3_51 in3_52 9.241569
Rin3_53 in3_52 in3_53 9.241569
Rin3_54 in3_53 in3_54 9.241569
Rin3_55 in3_54 in3_55 9.241569
Rin3_56 in3_55 in3_56 9.241569
Rin3_57 in3 in3_57 9.241569
Rin3_58 in3_57 in3_58 9.241569
Rin3_59 in3_58 in3_59 9.241569
Rin3_60 in3_59 in3_60 9.241569
Rin3_61 in3_60 in3_61 9.241569
Rin3_62 in3_61 in3_62 9.241569
Rin3_63 in3_62 in3_63 9.241569
Rin3_64 in3_63 in3_64 9.241569
Rin3_65 in3_64 in3_65 9.241569
Rin3_66 in3_65 in3_66 9.241569
Rin3_67 in3_66 in3_67 9.241569
Rin3_68 in3_67 in3_68 9.241569
Rin3_69 in3_68 in3_69 9.241569
Rin3_70 in3_69 in3_70 9.241569
Rin3_71 in3_70 in3_71 9.241569
Rin3_72 in3_71 in3_72 9.241569
Rin3_73 in3_72 in3_73 9.241569
Rin3_74 in3_73 in3_74 9.241569
Rin3_75 in3_74 in3_75 9.241569
Rin3_76 in3_75 in3_76 9.241569
Rin3_77 in3_76 in3_77 9.241569
Rin3_78 in3_77 in3_78 9.241569
Rin3_79 in3_78 in3_79 9.241569
Rin3_80 in3_79 in3_80 9.241569
Rin3_81 in3_80 in3_81 9.241569
Rin3_82 in3_81 in3_82 9.241569
Rin3_83 in3_82 in3_83 9.241569
Rin3_84 in3_83 in3_84 9.241569
Rin4_1 in4 in4_1 9.241569
Rin4_2 in4_1 in4_2 9.241569
Rin4_3 in4_2 in4_3 9.241569
Rin4_4 in4_3 in4_4 9.241569
Rin4_5 in4_4 in4_5 9.241569
Rin4_6 in4_5 in4_6 9.241569
Rin4_7 in4_6 in4_7 9.241569
Rin4_8 in4_7 in4_8 9.241569
Rin4_9 in4_8 in4_9 9.241569
Rin4_10 in4_9 in4_10 9.241569
Rin4_11 in4_10 in4_11 9.241569
Rin4_12 in4_11 in4_12 9.241569
Rin4_13 in4_12 in4_13 9.241569
Rin4_14 in4_13 in4_14 9.241569
Rin4_15 in4_14 in4_15 9.241569
Rin4_16 in4_15 in4_16 9.241569
Rin4_17 in4_16 in4_17 9.241569
Rin4_18 in4_17 in4_18 9.241569
Rin4_19 in4_18 in4_19 9.241569
Rin4_20 in4_19 in4_20 9.241569
Rin4_21 in4_20 in4_21 9.241569
Rin4_22 in4_21 in4_22 9.241569
Rin4_23 in4_22 in4_23 9.241569
Rin4_24 in4_23 in4_24 9.241569
Rin4_25 in4_24 in4_25 9.241569
Rin4_26 in4_25 in4_26 9.241569
Rin4_27 in4_26 in4_27 9.241569
Rin4_28 in4_27 in4_28 9.241569
Rin4_29 in4 in4_29 9.241569
Rin4_30 in4_29 in4_30 9.241569
Rin4_31 in4_30 in4_31 9.241569
Rin4_32 in4_31 in4_32 9.241569
Rin4_33 in4_32 in4_33 9.241569
Rin4_34 in4_33 in4_34 9.241569
Rin4_35 in4_34 in4_35 9.241569
Rin4_36 in4_35 in4_36 9.241569
Rin4_37 in4_36 in4_37 9.241569
Rin4_38 in4_37 in4_38 9.241569
Rin4_39 in4_38 in4_39 9.241569
Rin4_40 in4_39 in4_40 9.241569
Rin4_41 in4_40 in4_41 9.241569
Rin4_42 in4_41 in4_42 9.241569
Rin4_43 in4_42 in4_43 9.241569
Rin4_44 in4_43 in4_44 9.241569
Rin4_45 in4_44 in4_45 9.241569
Rin4_46 in4_45 in4_46 9.241569
Rin4_47 in4_46 in4_47 9.241569
Rin4_48 in4_47 in4_48 9.241569
Rin4_49 in4_48 in4_49 9.241569
Rin4_50 in4_49 in4_50 9.241569
Rin4_51 in4_50 in4_51 9.241569
Rin4_52 in4_51 in4_52 9.241569
Rin4_53 in4_52 in4_53 9.241569
Rin4_54 in4_53 in4_54 9.241569
Rin4_55 in4_54 in4_55 9.241569
Rin4_56 in4_55 in4_56 9.241569
Rin4_57 in4 in4_57 9.241569
Rin4_58 in4_57 in4_58 9.241569
Rin4_59 in4_58 in4_59 9.241569
Rin4_60 in4_59 in4_60 9.241569
Rin4_61 in4_60 in4_61 9.241569
Rin4_62 in4_61 in4_62 9.241569
Rin4_63 in4_62 in4_63 9.241569
Rin4_64 in4_63 in4_64 9.241569
Rin4_65 in4_64 in4_65 9.241569
Rin4_66 in4_65 in4_66 9.241569
Rin4_67 in4_66 in4_67 9.241569
Rin4_68 in4_67 in4_68 9.241569
Rin4_69 in4_68 in4_69 9.241569
Rin4_70 in4_69 in4_70 9.241569
Rin4_71 in4_70 in4_71 9.241569
Rin4_72 in4_71 in4_72 9.241569
Rin4_73 in4_72 in4_73 9.241569
Rin4_74 in4_73 in4_74 9.241569
Rin4_75 in4_74 in4_75 9.241569
Rin4_76 in4_75 in4_76 9.241569
Rin4_77 in4_76 in4_77 9.241569
Rin4_78 in4_77 in4_78 9.241569
Rin4_79 in4_78 in4_79 9.241569
Rin4_80 in4_79 in4_80 9.241569
Rin4_81 in4_80 in4_81 9.241569
Rin4_82 in4_81 in4_82 9.241569
Rin4_83 in4_82 in4_83 9.241569
Rin4_84 in4_83 in4_84 9.241569
Rin5_1 in5 in5_1 9.241569
Rin5_2 in5_1 in5_2 9.241569
Rin5_3 in5_2 in5_3 9.241569
Rin5_4 in5_3 in5_4 9.241569
Rin5_5 in5_4 in5_5 9.241569
Rin5_6 in5_5 in5_6 9.241569
Rin5_7 in5_6 in5_7 9.241569
Rin5_8 in5_7 in5_8 9.241569
Rin5_9 in5_8 in5_9 9.241569
Rin5_10 in5_9 in5_10 9.241569
Rin5_11 in5_10 in5_11 9.241569
Rin5_12 in5_11 in5_12 9.241569
Rin5_13 in5_12 in5_13 9.241569
Rin5_14 in5_13 in5_14 9.241569
Rin5_15 in5_14 in5_15 9.241569
Rin5_16 in5_15 in5_16 9.241569
Rin5_17 in5_16 in5_17 9.241569
Rin5_18 in5_17 in5_18 9.241569
Rin5_19 in5_18 in5_19 9.241569
Rin5_20 in5_19 in5_20 9.241569
Rin5_21 in5_20 in5_21 9.241569
Rin5_22 in5_21 in5_22 9.241569
Rin5_23 in5_22 in5_23 9.241569
Rin5_24 in5_23 in5_24 9.241569
Rin5_25 in5_24 in5_25 9.241569
Rin5_26 in5_25 in5_26 9.241569
Rin5_27 in5_26 in5_27 9.241569
Rin5_28 in5_27 in5_28 9.241569
Rin5_29 in5 in5_29 9.241569
Rin5_30 in5_29 in5_30 9.241569
Rin5_31 in5_30 in5_31 9.241569
Rin5_32 in5_31 in5_32 9.241569
Rin5_33 in5_32 in5_33 9.241569
Rin5_34 in5_33 in5_34 9.241569
Rin5_35 in5_34 in5_35 9.241569
Rin5_36 in5_35 in5_36 9.241569
Rin5_37 in5_36 in5_37 9.241569
Rin5_38 in5_37 in5_38 9.241569
Rin5_39 in5_38 in5_39 9.241569
Rin5_40 in5_39 in5_40 9.241569
Rin5_41 in5_40 in5_41 9.241569
Rin5_42 in5_41 in5_42 9.241569
Rin5_43 in5_42 in5_43 9.241569
Rin5_44 in5_43 in5_44 9.241569
Rin5_45 in5_44 in5_45 9.241569
Rin5_46 in5_45 in5_46 9.241569
Rin5_47 in5_46 in5_47 9.241569
Rin5_48 in5_47 in5_48 9.241569
Rin5_49 in5_48 in5_49 9.241569
Rin5_50 in5_49 in5_50 9.241569
Rin5_51 in5_50 in5_51 9.241569
Rin5_52 in5_51 in5_52 9.241569
Rin5_53 in5_52 in5_53 9.241569
Rin5_54 in5_53 in5_54 9.241569
Rin5_55 in5_54 in5_55 9.241569
Rin5_56 in5_55 in5_56 9.241569
Rin5_57 in5 in5_57 9.241569
Rin5_58 in5_57 in5_58 9.241569
Rin5_59 in5_58 in5_59 9.241569
Rin5_60 in5_59 in5_60 9.241569
Rin5_61 in5_60 in5_61 9.241569
Rin5_62 in5_61 in5_62 9.241569
Rin5_63 in5_62 in5_63 9.241569
Rin5_64 in5_63 in5_64 9.241569
Rin5_65 in5_64 in5_65 9.241569
Rin5_66 in5_65 in5_66 9.241569
Rin5_67 in5_66 in5_67 9.241569
Rin5_68 in5_67 in5_68 9.241569
Rin5_69 in5_68 in5_69 9.241569
Rin5_70 in5_69 in5_70 9.241569
Rin5_71 in5_70 in5_71 9.241569
Rin5_72 in5_71 in5_72 9.241569
Rin5_73 in5_72 in5_73 9.241569
Rin5_74 in5_73 in5_74 9.241569
Rin5_75 in5_74 in5_75 9.241569
Rin5_76 in5_75 in5_76 9.241569
Rin5_77 in5_76 in5_77 9.241569
Rin5_78 in5_77 in5_78 9.241569
Rin5_79 in5_78 in5_79 9.241569
Rin5_80 in5_79 in5_80 9.241569
Rin5_81 in5_80 in5_81 9.241569
Rin5_82 in5_81 in5_82 9.241569
Rin5_83 in5_82 in5_83 9.241569
Rin5_84 in5_83 in5_84 9.241569
Rin6_1 in6 in6_1 9.241569
Rin6_2 in6_1 in6_2 9.241569
Rin6_3 in6_2 in6_3 9.241569
Rin6_4 in6_3 in6_4 9.241569
Rin6_5 in6_4 in6_5 9.241569
Rin6_6 in6_5 in6_6 9.241569
Rin6_7 in6_6 in6_7 9.241569
Rin6_8 in6_7 in6_8 9.241569
Rin6_9 in6_8 in6_9 9.241569
Rin6_10 in6_9 in6_10 9.241569
Rin6_11 in6_10 in6_11 9.241569
Rin6_12 in6_11 in6_12 9.241569
Rin6_13 in6_12 in6_13 9.241569
Rin6_14 in6_13 in6_14 9.241569
Rin6_15 in6_14 in6_15 9.241569
Rin6_16 in6_15 in6_16 9.241569
Rin6_17 in6_16 in6_17 9.241569
Rin6_18 in6_17 in6_18 9.241569
Rin6_19 in6_18 in6_19 9.241569
Rin6_20 in6_19 in6_20 9.241569
Rin6_21 in6_20 in6_21 9.241569
Rin6_22 in6_21 in6_22 9.241569
Rin6_23 in6_22 in6_23 9.241569
Rin6_24 in6_23 in6_24 9.241569
Rin6_25 in6_24 in6_25 9.241569
Rin6_26 in6_25 in6_26 9.241569
Rin6_27 in6_26 in6_27 9.241569
Rin6_28 in6_27 in6_28 9.241569
Rin6_29 in6 in6_29 9.241569
Rin6_30 in6_29 in6_30 9.241569
Rin6_31 in6_30 in6_31 9.241569
Rin6_32 in6_31 in6_32 9.241569
Rin6_33 in6_32 in6_33 9.241569
Rin6_34 in6_33 in6_34 9.241569
Rin6_35 in6_34 in6_35 9.241569
Rin6_36 in6_35 in6_36 9.241569
Rin6_37 in6_36 in6_37 9.241569
Rin6_38 in6_37 in6_38 9.241569
Rin6_39 in6_38 in6_39 9.241569
Rin6_40 in6_39 in6_40 9.241569
Rin6_41 in6_40 in6_41 9.241569
Rin6_42 in6_41 in6_42 9.241569
Rin6_43 in6_42 in6_43 9.241569
Rin6_44 in6_43 in6_44 9.241569
Rin6_45 in6_44 in6_45 9.241569
Rin6_46 in6_45 in6_46 9.241569
Rin6_47 in6_46 in6_47 9.241569
Rin6_48 in6_47 in6_48 9.241569
Rin6_49 in6_48 in6_49 9.241569
Rin6_50 in6_49 in6_50 9.241569
Rin6_51 in6_50 in6_51 9.241569
Rin6_52 in6_51 in6_52 9.241569
Rin6_53 in6_52 in6_53 9.241569
Rin6_54 in6_53 in6_54 9.241569
Rin6_55 in6_54 in6_55 9.241569
Rin6_56 in6_55 in6_56 9.241569
Rin6_57 in6 in6_57 9.241569
Rin6_58 in6_57 in6_58 9.241569
Rin6_59 in6_58 in6_59 9.241569
Rin6_60 in6_59 in6_60 9.241569
Rin6_61 in6_60 in6_61 9.241569
Rin6_62 in6_61 in6_62 9.241569
Rin6_63 in6_62 in6_63 9.241569
Rin6_64 in6_63 in6_64 9.241569
Rin6_65 in6_64 in6_65 9.241569
Rin6_66 in6_65 in6_66 9.241569
Rin6_67 in6_66 in6_67 9.241569
Rin6_68 in6_67 in6_68 9.241569
Rin6_69 in6_68 in6_69 9.241569
Rin6_70 in6_69 in6_70 9.241569
Rin6_71 in6_70 in6_71 9.241569
Rin6_72 in6_71 in6_72 9.241569
Rin6_73 in6_72 in6_73 9.241569
Rin6_74 in6_73 in6_74 9.241569
Rin6_75 in6_74 in6_75 9.241569
Rin6_76 in6_75 in6_76 9.241569
Rin6_77 in6_76 in6_77 9.241569
Rin6_78 in6_77 in6_78 9.241569
Rin6_79 in6_78 in6_79 9.241569
Rin6_80 in6_79 in6_80 9.241569
Rin6_81 in6_80 in6_81 9.241569
Rin6_82 in6_81 in6_82 9.241569
Rin6_83 in6_82 in6_83 9.241569
Rin6_84 in6_83 in6_84 9.241569
Rin7_1 in7 in7_1 9.241569
Rin7_2 in7_1 in7_2 9.241569
Rin7_3 in7_2 in7_3 9.241569
Rin7_4 in7_3 in7_4 9.241569
Rin7_5 in7_4 in7_5 9.241569
Rin7_6 in7_5 in7_6 9.241569
Rin7_7 in7_6 in7_7 9.241569
Rin7_8 in7_7 in7_8 9.241569
Rin7_9 in7_8 in7_9 9.241569
Rin7_10 in7_9 in7_10 9.241569
Rin7_11 in7_10 in7_11 9.241569
Rin7_12 in7_11 in7_12 9.241569
Rin7_13 in7_12 in7_13 9.241569
Rin7_14 in7_13 in7_14 9.241569
Rin7_15 in7_14 in7_15 9.241569
Rin7_16 in7_15 in7_16 9.241569
Rin7_17 in7_16 in7_17 9.241569
Rin7_18 in7_17 in7_18 9.241569
Rin7_19 in7_18 in7_19 9.241569
Rin7_20 in7_19 in7_20 9.241569
Rin7_21 in7_20 in7_21 9.241569
Rin7_22 in7_21 in7_22 9.241569
Rin7_23 in7_22 in7_23 9.241569
Rin7_24 in7_23 in7_24 9.241569
Rin7_25 in7_24 in7_25 9.241569
Rin7_26 in7_25 in7_26 9.241569
Rin7_27 in7_26 in7_27 9.241569
Rin7_28 in7_27 in7_28 9.241569
Rin7_29 in7 in7_29 9.241569
Rin7_30 in7_29 in7_30 9.241569
Rin7_31 in7_30 in7_31 9.241569
Rin7_32 in7_31 in7_32 9.241569
Rin7_33 in7_32 in7_33 9.241569
Rin7_34 in7_33 in7_34 9.241569
Rin7_35 in7_34 in7_35 9.241569
Rin7_36 in7_35 in7_36 9.241569
Rin7_37 in7_36 in7_37 9.241569
Rin7_38 in7_37 in7_38 9.241569
Rin7_39 in7_38 in7_39 9.241569
Rin7_40 in7_39 in7_40 9.241569
Rin7_41 in7_40 in7_41 9.241569
Rin7_42 in7_41 in7_42 9.241569
Rin7_43 in7_42 in7_43 9.241569
Rin7_44 in7_43 in7_44 9.241569
Rin7_45 in7_44 in7_45 9.241569
Rin7_46 in7_45 in7_46 9.241569
Rin7_47 in7_46 in7_47 9.241569
Rin7_48 in7_47 in7_48 9.241569
Rin7_49 in7_48 in7_49 9.241569
Rin7_50 in7_49 in7_50 9.241569
Rin7_51 in7_50 in7_51 9.241569
Rin7_52 in7_51 in7_52 9.241569
Rin7_53 in7_52 in7_53 9.241569
Rin7_54 in7_53 in7_54 9.241569
Rin7_55 in7_54 in7_55 9.241569
Rin7_56 in7_55 in7_56 9.241569
Rin7_57 in7 in7_57 9.241569
Rin7_58 in7_57 in7_58 9.241569
Rin7_59 in7_58 in7_59 9.241569
Rin7_60 in7_59 in7_60 9.241569
Rin7_61 in7_60 in7_61 9.241569
Rin7_62 in7_61 in7_62 9.241569
Rin7_63 in7_62 in7_63 9.241569
Rin7_64 in7_63 in7_64 9.241569
Rin7_65 in7_64 in7_65 9.241569
Rin7_66 in7_65 in7_66 9.241569
Rin7_67 in7_66 in7_67 9.241569
Rin7_68 in7_67 in7_68 9.241569
Rin7_69 in7_68 in7_69 9.241569
Rin7_70 in7_69 in7_70 9.241569
Rin7_71 in7_70 in7_71 9.241569
Rin7_72 in7_71 in7_72 9.241569
Rin7_73 in7_72 in7_73 9.241569
Rin7_74 in7_73 in7_74 9.241569
Rin7_75 in7_74 in7_75 9.241569
Rin7_76 in7_75 in7_76 9.241569
Rin7_77 in7_76 in7_77 9.241569
Rin7_78 in7_77 in7_78 9.241569
Rin7_79 in7_78 in7_79 9.241569
Rin7_80 in7_79 in7_80 9.241569
Rin7_81 in7_80 in7_81 9.241569
Rin7_82 in7_81 in7_82 9.241569
Rin7_83 in7_82 in7_83 9.241569
Rin7_84 in7_83 in7_84 9.241569
Rin8_1 in8 in8_1 9.241569
Rin8_2 in8_1 in8_2 9.241569
Rin8_3 in8_2 in8_3 9.241569
Rin8_4 in8_3 in8_4 9.241569
Rin8_5 in8_4 in8_5 9.241569
Rin8_6 in8_5 in8_6 9.241569
Rin8_7 in8_6 in8_7 9.241569
Rin8_8 in8_7 in8_8 9.241569
Rin8_9 in8_8 in8_9 9.241569
Rin8_10 in8_9 in8_10 9.241569
Rin8_11 in8_10 in8_11 9.241569
Rin8_12 in8_11 in8_12 9.241569
Rin8_13 in8_12 in8_13 9.241569
Rin8_14 in8_13 in8_14 9.241569
Rin8_15 in8_14 in8_15 9.241569
Rin8_16 in8_15 in8_16 9.241569
Rin8_17 in8_16 in8_17 9.241569
Rin8_18 in8_17 in8_18 9.241569
Rin8_19 in8_18 in8_19 9.241569
Rin8_20 in8_19 in8_20 9.241569
Rin8_21 in8_20 in8_21 9.241569
Rin8_22 in8_21 in8_22 9.241569
Rin8_23 in8_22 in8_23 9.241569
Rin8_24 in8_23 in8_24 9.241569
Rin8_25 in8_24 in8_25 9.241569
Rin8_26 in8_25 in8_26 9.241569
Rin8_27 in8_26 in8_27 9.241569
Rin8_28 in8_27 in8_28 9.241569
Rin8_29 in8 in8_29 9.241569
Rin8_30 in8_29 in8_30 9.241569
Rin8_31 in8_30 in8_31 9.241569
Rin8_32 in8_31 in8_32 9.241569
Rin8_33 in8_32 in8_33 9.241569
Rin8_34 in8_33 in8_34 9.241569
Rin8_35 in8_34 in8_35 9.241569
Rin8_36 in8_35 in8_36 9.241569
Rin8_37 in8_36 in8_37 9.241569
Rin8_38 in8_37 in8_38 9.241569
Rin8_39 in8_38 in8_39 9.241569
Rin8_40 in8_39 in8_40 9.241569
Rin8_41 in8_40 in8_41 9.241569
Rin8_42 in8_41 in8_42 9.241569
Rin8_43 in8_42 in8_43 9.241569
Rin8_44 in8_43 in8_44 9.241569
Rin8_45 in8_44 in8_45 9.241569
Rin8_46 in8_45 in8_46 9.241569
Rin8_47 in8_46 in8_47 9.241569
Rin8_48 in8_47 in8_48 9.241569
Rin8_49 in8_48 in8_49 9.241569
Rin8_50 in8_49 in8_50 9.241569
Rin8_51 in8_50 in8_51 9.241569
Rin8_52 in8_51 in8_52 9.241569
Rin8_53 in8_52 in8_53 9.241569
Rin8_54 in8_53 in8_54 9.241569
Rin8_55 in8_54 in8_55 9.241569
Rin8_56 in8_55 in8_56 9.241569
Rin8_57 in8 in8_57 9.241569
Rin8_58 in8_57 in8_58 9.241569
Rin8_59 in8_58 in8_59 9.241569
Rin8_60 in8_59 in8_60 9.241569
Rin8_61 in8_60 in8_61 9.241569
Rin8_62 in8_61 in8_62 9.241569
Rin8_63 in8_62 in8_63 9.241569
Rin8_64 in8_63 in8_64 9.241569
Rin8_65 in8_64 in8_65 9.241569
Rin8_66 in8_65 in8_66 9.241569
Rin8_67 in8_66 in8_67 9.241569
Rin8_68 in8_67 in8_68 9.241569
Rin8_69 in8_68 in8_69 9.241569
Rin8_70 in8_69 in8_70 9.241569
Rin8_71 in8_70 in8_71 9.241569
Rin8_72 in8_71 in8_72 9.241569
Rin8_73 in8_72 in8_73 9.241569
Rin8_74 in8_73 in8_74 9.241569
Rin8_75 in8_74 in8_75 9.241569
Rin8_76 in8_75 in8_76 9.241569
Rin8_77 in8_76 in8_77 9.241569
Rin8_78 in8_77 in8_78 9.241569
Rin8_79 in8_78 in8_79 9.241569
Rin8_80 in8_79 in8_80 9.241569
Rin8_81 in8_80 in8_81 9.241569
Rin8_82 in8_81 in8_82 9.241569
Rin8_83 in8_82 in8_83 9.241569
Rin8_84 in8_83 in8_84 9.241569
Rin9_1 in9 in9_1 9.241569
Rin9_2 in9_1 in9_2 9.241569
Rin9_3 in9_2 in9_3 9.241569
Rin9_4 in9_3 in9_4 9.241569
Rin9_5 in9_4 in9_5 9.241569
Rin9_6 in9_5 in9_6 9.241569
Rin9_7 in9_6 in9_7 9.241569
Rin9_8 in9_7 in9_8 9.241569
Rin9_9 in9_8 in9_9 9.241569
Rin9_10 in9_9 in9_10 9.241569
Rin9_11 in9_10 in9_11 9.241569
Rin9_12 in9_11 in9_12 9.241569
Rin9_13 in9_12 in9_13 9.241569
Rin9_14 in9_13 in9_14 9.241569
Rin9_15 in9_14 in9_15 9.241569
Rin9_16 in9_15 in9_16 9.241569
Rin9_17 in9_16 in9_17 9.241569
Rin9_18 in9_17 in9_18 9.241569
Rin9_19 in9_18 in9_19 9.241569
Rin9_20 in9_19 in9_20 9.241569
Rin9_21 in9_20 in9_21 9.241569
Rin9_22 in9_21 in9_22 9.241569
Rin9_23 in9_22 in9_23 9.241569
Rin9_24 in9_23 in9_24 9.241569
Rin9_25 in9_24 in9_25 9.241569
Rin9_26 in9_25 in9_26 9.241569
Rin9_27 in9_26 in9_27 9.241569
Rin9_28 in9_27 in9_28 9.241569
Rin9_29 in9 in9_29 9.241569
Rin9_30 in9_29 in9_30 9.241569
Rin9_31 in9_30 in9_31 9.241569
Rin9_32 in9_31 in9_32 9.241569
Rin9_33 in9_32 in9_33 9.241569
Rin9_34 in9_33 in9_34 9.241569
Rin9_35 in9_34 in9_35 9.241569
Rin9_36 in9_35 in9_36 9.241569
Rin9_37 in9_36 in9_37 9.241569
Rin9_38 in9_37 in9_38 9.241569
Rin9_39 in9_38 in9_39 9.241569
Rin9_40 in9_39 in9_40 9.241569
Rin9_41 in9_40 in9_41 9.241569
Rin9_42 in9_41 in9_42 9.241569
Rin9_43 in9_42 in9_43 9.241569
Rin9_44 in9_43 in9_44 9.241569
Rin9_45 in9_44 in9_45 9.241569
Rin9_46 in9_45 in9_46 9.241569
Rin9_47 in9_46 in9_47 9.241569
Rin9_48 in9_47 in9_48 9.241569
Rin9_49 in9_48 in9_49 9.241569
Rin9_50 in9_49 in9_50 9.241569
Rin9_51 in9_50 in9_51 9.241569
Rin9_52 in9_51 in9_52 9.241569
Rin9_53 in9_52 in9_53 9.241569
Rin9_54 in9_53 in9_54 9.241569
Rin9_55 in9_54 in9_55 9.241569
Rin9_56 in9_55 in9_56 9.241569
Rin9_57 in9 in9_57 9.241569
Rin9_58 in9_57 in9_58 9.241569
Rin9_59 in9_58 in9_59 9.241569
Rin9_60 in9_59 in9_60 9.241569
Rin9_61 in9_60 in9_61 9.241569
Rin9_62 in9_61 in9_62 9.241569
Rin9_63 in9_62 in9_63 9.241569
Rin9_64 in9_63 in9_64 9.241569
Rin9_65 in9_64 in9_65 9.241569
Rin9_66 in9_65 in9_66 9.241569
Rin9_67 in9_66 in9_67 9.241569
Rin9_68 in9_67 in9_68 9.241569
Rin9_69 in9_68 in9_69 9.241569
Rin9_70 in9_69 in9_70 9.241569
Rin9_71 in9_70 in9_71 9.241569
Rin9_72 in9_71 in9_72 9.241569
Rin9_73 in9_72 in9_73 9.241569
Rin9_74 in9_73 in9_74 9.241569
Rin9_75 in9_74 in9_75 9.241569
Rin9_76 in9_75 in9_76 9.241569
Rin9_77 in9_76 in9_77 9.241569
Rin9_78 in9_77 in9_78 9.241569
Rin9_79 in9_78 in9_79 9.241569
Rin9_80 in9_79 in9_80 9.241569
Rin9_81 in9_80 in9_81 9.241569
Rin9_82 in9_81 in9_82 9.241569
Rin9_83 in9_82 in9_83 9.241569
Rin9_84 in9_83 in9_84 9.241569
Rin10_1 in10 in10_1 9.241569
Rin10_2 in10_1 in10_2 9.241569
Rin10_3 in10_2 in10_3 9.241569
Rin10_4 in10_3 in10_4 9.241569
Rin10_5 in10_4 in10_5 9.241569
Rin10_6 in10_5 in10_6 9.241569
Rin10_7 in10_6 in10_7 9.241569
Rin10_8 in10_7 in10_8 9.241569
Rin10_9 in10_8 in10_9 9.241569
Rin10_10 in10_9 in10_10 9.241569
Rin10_11 in10_10 in10_11 9.241569
Rin10_12 in10_11 in10_12 9.241569
Rin10_13 in10_12 in10_13 9.241569
Rin10_14 in10_13 in10_14 9.241569
Rin10_15 in10_14 in10_15 9.241569
Rin10_16 in10_15 in10_16 9.241569
Rin10_17 in10_16 in10_17 9.241569
Rin10_18 in10_17 in10_18 9.241569
Rin10_19 in10_18 in10_19 9.241569
Rin10_20 in10_19 in10_20 9.241569
Rin10_21 in10_20 in10_21 9.241569
Rin10_22 in10_21 in10_22 9.241569
Rin10_23 in10_22 in10_23 9.241569
Rin10_24 in10_23 in10_24 9.241569
Rin10_25 in10_24 in10_25 9.241569
Rin10_26 in10_25 in10_26 9.241569
Rin10_27 in10_26 in10_27 9.241569
Rin10_28 in10_27 in10_28 9.241569
Rin10_29 in10 in10_29 9.241569
Rin10_30 in10_29 in10_30 9.241569
Rin10_31 in10_30 in10_31 9.241569
Rin10_32 in10_31 in10_32 9.241569
Rin10_33 in10_32 in10_33 9.241569
Rin10_34 in10_33 in10_34 9.241569
Rin10_35 in10_34 in10_35 9.241569
Rin10_36 in10_35 in10_36 9.241569
Rin10_37 in10_36 in10_37 9.241569
Rin10_38 in10_37 in10_38 9.241569
Rin10_39 in10_38 in10_39 9.241569
Rin10_40 in10_39 in10_40 9.241569
Rin10_41 in10_40 in10_41 9.241569
Rin10_42 in10_41 in10_42 9.241569
Rin10_43 in10_42 in10_43 9.241569
Rin10_44 in10_43 in10_44 9.241569
Rin10_45 in10_44 in10_45 9.241569
Rin10_46 in10_45 in10_46 9.241569
Rin10_47 in10_46 in10_47 9.241569
Rin10_48 in10_47 in10_48 9.241569
Rin10_49 in10_48 in10_49 9.241569
Rin10_50 in10_49 in10_50 9.241569
Rin10_51 in10_50 in10_51 9.241569
Rin10_52 in10_51 in10_52 9.241569
Rin10_53 in10_52 in10_53 9.241569
Rin10_54 in10_53 in10_54 9.241569
Rin10_55 in10_54 in10_55 9.241569
Rin10_56 in10_55 in10_56 9.241569
Rin10_57 in10 in10_57 9.241569
Rin10_58 in10_57 in10_58 9.241569
Rin10_59 in10_58 in10_59 9.241569
Rin10_60 in10_59 in10_60 9.241569
Rin10_61 in10_60 in10_61 9.241569
Rin10_62 in10_61 in10_62 9.241569
Rin10_63 in10_62 in10_63 9.241569
Rin10_64 in10_63 in10_64 9.241569
Rin10_65 in10_64 in10_65 9.241569
Rin10_66 in10_65 in10_66 9.241569
Rin10_67 in10_66 in10_67 9.241569
Rin10_68 in10_67 in10_68 9.241569
Rin10_69 in10_68 in10_69 9.241569
Rin10_70 in10_69 in10_70 9.241569
Rin10_71 in10_70 in10_71 9.241569
Rin10_72 in10_71 in10_72 9.241569
Rin10_73 in10_72 in10_73 9.241569
Rin10_74 in10_73 in10_74 9.241569
Rin10_75 in10_74 in10_75 9.241569
Rin10_76 in10_75 in10_76 9.241569
Rin10_77 in10_76 in10_77 9.241569
Rin10_78 in10_77 in10_78 9.241569
Rin10_79 in10_78 in10_79 9.241569
Rin10_80 in10_79 in10_80 9.241569
Rin10_81 in10_80 in10_81 9.241569
Rin10_82 in10_81 in10_82 9.241569
Rin10_83 in10_82 in10_83 9.241569
Rin10_84 in10_83 in10_84 9.241569
Rin11_1 in11 in11_1 9.241569
Rin11_2 in11_1 in11_2 9.241569
Rin11_3 in11_2 in11_3 9.241569
Rin11_4 in11_3 in11_4 9.241569
Rin11_5 in11_4 in11_5 9.241569
Rin11_6 in11_5 in11_6 9.241569
Rin11_7 in11_6 in11_7 9.241569
Rin11_8 in11_7 in11_8 9.241569
Rin11_9 in11_8 in11_9 9.241569
Rin11_10 in11_9 in11_10 9.241569
Rin11_11 in11_10 in11_11 9.241569
Rin11_12 in11_11 in11_12 9.241569
Rin11_13 in11_12 in11_13 9.241569
Rin11_14 in11_13 in11_14 9.241569
Rin11_15 in11_14 in11_15 9.241569
Rin11_16 in11_15 in11_16 9.241569
Rin11_17 in11_16 in11_17 9.241569
Rin11_18 in11_17 in11_18 9.241569
Rin11_19 in11_18 in11_19 9.241569
Rin11_20 in11_19 in11_20 9.241569
Rin11_21 in11_20 in11_21 9.241569
Rin11_22 in11_21 in11_22 9.241569
Rin11_23 in11_22 in11_23 9.241569
Rin11_24 in11_23 in11_24 9.241569
Rin11_25 in11_24 in11_25 9.241569
Rin11_26 in11_25 in11_26 9.241569
Rin11_27 in11_26 in11_27 9.241569
Rin11_28 in11_27 in11_28 9.241569
Rin11_29 in11 in11_29 9.241569
Rin11_30 in11_29 in11_30 9.241569
Rin11_31 in11_30 in11_31 9.241569
Rin11_32 in11_31 in11_32 9.241569
Rin11_33 in11_32 in11_33 9.241569
Rin11_34 in11_33 in11_34 9.241569
Rin11_35 in11_34 in11_35 9.241569
Rin11_36 in11_35 in11_36 9.241569
Rin11_37 in11_36 in11_37 9.241569
Rin11_38 in11_37 in11_38 9.241569
Rin11_39 in11_38 in11_39 9.241569
Rin11_40 in11_39 in11_40 9.241569
Rin11_41 in11_40 in11_41 9.241569
Rin11_42 in11_41 in11_42 9.241569
Rin11_43 in11_42 in11_43 9.241569
Rin11_44 in11_43 in11_44 9.241569
Rin11_45 in11_44 in11_45 9.241569
Rin11_46 in11_45 in11_46 9.241569
Rin11_47 in11_46 in11_47 9.241569
Rin11_48 in11_47 in11_48 9.241569
Rin11_49 in11_48 in11_49 9.241569
Rin11_50 in11_49 in11_50 9.241569
Rin11_51 in11_50 in11_51 9.241569
Rin11_52 in11_51 in11_52 9.241569
Rin11_53 in11_52 in11_53 9.241569
Rin11_54 in11_53 in11_54 9.241569
Rin11_55 in11_54 in11_55 9.241569
Rin11_56 in11_55 in11_56 9.241569
Rin11_57 in11 in11_57 9.241569
Rin11_58 in11_57 in11_58 9.241569
Rin11_59 in11_58 in11_59 9.241569
Rin11_60 in11_59 in11_60 9.241569
Rin11_61 in11_60 in11_61 9.241569
Rin11_62 in11_61 in11_62 9.241569
Rin11_63 in11_62 in11_63 9.241569
Rin11_64 in11_63 in11_64 9.241569
Rin11_65 in11_64 in11_65 9.241569
Rin11_66 in11_65 in11_66 9.241569
Rin11_67 in11_66 in11_67 9.241569
Rin11_68 in11_67 in11_68 9.241569
Rin11_69 in11_68 in11_69 9.241569
Rin11_70 in11_69 in11_70 9.241569
Rin11_71 in11_70 in11_71 9.241569
Rin11_72 in11_71 in11_72 9.241569
Rin11_73 in11_72 in11_73 9.241569
Rin11_74 in11_73 in11_74 9.241569
Rin11_75 in11_74 in11_75 9.241569
Rin11_76 in11_75 in11_76 9.241569
Rin11_77 in11_76 in11_77 9.241569
Rin11_78 in11_77 in11_78 9.241569
Rin11_79 in11_78 in11_79 9.241569
Rin11_80 in11_79 in11_80 9.241569
Rin11_81 in11_80 in11_81 9.241569
Rin11_82 in11_81 in11_82 9.241569
Rin11_83 in11_82 in11_83 9.241569
Rin11_84 in11_83 in11_84 9.241569
Rin12_1 in12 in12_1 9.241569
Rin12_2 in12_1 in12_2 9.241569
Rin12_3 in12_2 in12_3 9.241569
Rin12_4 in12_3 in12_4 9.241569
Rin12_5 in12_4 in12_5 9.241569
Rin12_6 in12_5 in12_6 9.241569
Rin12_7 in12_6 in12_7 9.241569
Rin12_8 in12_7 in12_8 9.241569
Rin12_9 in12_8 in12_9 9.241569
Rin12_10 in12_9 in12_10 9.241569
Rin12_11 in12_10 in12_11 9.241569
Rin12_12 in12_11 in12_12 9.241569
Rin12_13 in12_12 in12_13 9.241569
Rin12_14 in12_13 in12_14 9.241569
Rin12_15 in12_14 in12_15 9.241569
Rin12_16 in12_15 in12_16 9.241569
Rin12_17 in12_16 in12_17 9.241569
Rin12_18 in12_17 in12_18 9.241569
Rin12_19 in12_18 in12_19 9.241569
Rin12_20 in12_19 in12_20 9.241569
Rin12_21 in12_20 in12_21 9.241569
Rin12_22 in12_21 in12_22 9.241569
Rin12_23 in12_22 in12_23 9.241569
Rin12_24 in12_23 in12_24 9.241569
Rin12_25 in12_24 in12_25 9.241569
Rin12_26 in12_25 in12_26 9.241569
Rin12_27 in12_26 in12_27 9.241569
Rin12_28 in12_27 in12_28 9.241569
Rin12_29 in12 in12_29 9.241569
Rin12_30 in12_29 in12_30 9.241569
Rin12_31 in12_30 in12_31 9.241569
Rin12_32 in12_31 in12_32 9.241569
Rin12_33 in12_32 in12_33 9.241569
Rin12_34 in12_33 in12_34 9.241569
Rin12_35 in12_34 in12_35 9.241569
Rin12_36 in12_35 in12_36 9.241569
Rin12_37 in12_36 in12_37 9.241569
Rin12_38 in12_37 in12_38 9.241569
Rin12_39 in12_38 in12_39 9.241569
Rin12_40 in12_39 in12_40 9.241569
Rin12_41 in12_40 in12_41 9.241569
Rin12_42 in12_41 in12_42 9.241569
Rin12_43 in12_42 in12_43 9.241569
Rin12_44 in12_43 in12_44 9.241569
Rin12_45 in12_44 in12_45 9.241569
Rin12_46 in12_45 in12_46 9.241569
Rin12_47 in12_46 in12_47 9.241569
Rin12_48 in12_47 in12_48 9.241569
Rin12_49 in12_48 in12_49 9.241569
Rin12_50 in12_49 in12_50 9.241569
Rin12_51 in12_50 in12_51 9.241569
Rin12_52 in12_51 in12_52 9.241569
Rin12_53 in12_52 in12_53 9.241569
Rin12_54 in12_53 in12_54 9.241569
Rin12_55 in12_54 in12_55 9.241569
Rin12_56 in12_55 in12_56 9.241569
Rin12_57 in12 in12_57 9.241569
Rin12_58 in12_57 in12_58 9.241569
Rin12_59 in12_58 in12_59 9.241569
Rin12_60 in12_59 in12_60 9.241569
Rin12_61 in12_60 in12_61 9.241569
Rin12_62 in12_61 in12_62 9.241569
Rin12_63 in12_62 in12_63 9.241569
Rin12_64 in12_63 in12_64 9.241569
Rin12_65 in12_64 in12_65 9.241569
Rin12_66 in12_65 in12_66 9.241569
Rin12_67 in12_66 in12_67 9.241569
Rin12_68 in12_67 in12_68 9.241569
Rin12_69 in12_68 in12_69 9.241569
Rin12_70 in12_69 in12_70 9.241569
Rin12_71 in12_70 in12_71 9.241569
Rin12_72 in12_71 in12_72 9.241569
Rin12_73 in12_72 in12_73 9.241569
Rin12_74 in12_73 in12_74 9.241569
Rin12_75 in12_74 in12_75 9.241569
Rin12_76 in12_75 in12_76 9.241569
Rin12_77 in12_76 in12_77 9.241569
Rin12_78 in12_77 in12_78 9.241569
Rin12_79 in12_78 in12_79 9.241569
Rin12_80 in12_79 in12_80 9.241569
Rin12_81 in12_80 in12_81 9.241569
Rin12_82 in12_81 in12_82 9.241569
Rin12_83 in12_82 in12_83 9.241569
Rin12_84 in12_83 in12_84 9.241569
Rin13_1 in13 in13_1 9.241569
Rin13_2 in13_1 in13_2 9.241569
Rin13_3 in13_2 in13_3 9.241569
Rin13_4 in13_3 in13_4 9.241569
Rin13_5 in13_4 in13_5 9.241569
Rin13_6 in13_5 in13_6 9.241569
Rin13_7 in13_6 in13_7 9.241569
Rin13_8 in13_7 in13_8 9.241569
Rin13_9 in13_8 in13_9 9.241569
Rin13_10 in13_9 in13_10 9.241569
Rin13_11 in13_10 in13_11 9.241569
Rin13_12 in13_11 in13_12 9.241569
Rin13_13 in13_12 in13_13 9.241569
Rin13_14 in13_13 in13_14 9.241569
Rin13_15 in13_14 in13_15 9.241569
Rin13_16 in13_15 in13_16 9.241569
Rin13_17 in13_16 in13_17 9.241569
Rin13_18 in13_17 in13_18 9.241569
Rin13_19 in13_18 in13_19 9.241569
Rin13_20 in13_19 in13_20 9.241569
Rin13_21 in13_20 in13_21 9.241569
Rin13_22 in13_21 in13_22 9.241569
Rin13_23 in13_22 in13_23 9.241569
Rin13_24 in13_23 in13_24 9.241569
Rin13_25 in13_24 in13_25 9.241569
Rin13_26 in13_25 in13_26 9.241569
Rin13_27 in13_26 in13_27 9.241569
Rin13_28 in13_27 in13_28 9.241569
Rin13_29 in13 in13_29 9.241569
Rin13_30 in13_29 in13_30 9.241569
Rin13_31 in13_30 in13_31 9.241569
Rin13_32 in13_31 in13_32 9.241569
Rin13_33 in13_32 in13_33 9.241569
Rin13_34 in13_33 in13_34 9.241569
Rin13_35 in13_34 in13_35 9.241569
Rin13_36 in13_35 in13_36 9.241569
Rin13_37 in13_36 in13_37 9.241569
Rin13_38 in13_37 in13_38 9.241569
Rin13_39 in13_38 in13_39 9.241569
Rin13_40 in13_39 in13_40 9.241569
Rin13_41 in13_40 in13_41 9.241569
Rin13_42 in13_41 in13_42 9.241569
Rin13_43 in13_42 in13_43 9.241569
Rin13_44 in13_43 in13_44 9.241569
Rin13_45 in13_44 in13_45 9.241569
Rin13_46 in13_45 in13_46 9.241569
Rin13_47 in13_46 in13_47 9.241569
Rin13_48 in13_47 in13_48 9.241569
Rin13_49 in13_48 in13_49 9.241569
Rin13_50 in13_49 in13_50 9.241569
Rin13_51 in13_50 in13_51 9.241569
Rin13_52 in13_51 in13_52 9.241569
Rin13_53 in13_52 in13_53 9.241569
Rin13_54 in13_53 in13_54 9.241569
Rin13_55 in13_54 in13_55 9.241569
Rin13_56 in13_55 in13_56 9.241569
Rin13_57 in13 in13_57 9.241569
Rin13_58 in13_57 in13_58 9.241569
Rin13_59 in13_58 in13_59 9.241569
Rin13_60 in13_59 in13_60 9.241569
Rin13_61 in13_60 in13_61 9.241569
Rin13_62 in13_61 in13_62 9.241569
Rin13_63 in13_62 in13_63 9.241569
Rin13_64 in13_63 in13_64 9.241569
Rin13_65 in13_64 in13_65 9.241569
Rin13_66 in13_65 in13_66 9.241569
Rin13_67 in13_66 in13_67 9.241569
Rin13_68 in13_67 in13_68 9.241569
Rin13_69 in13_68 in13_69 9.241569
Rin13_70 in13_69 in13_70 9.241569
Rin13_71 in13_70 in13_71 9.241569
Rin13_72 in13_71 in13_72 9.241569
Rin13_73 in13_72 in13_73 9.241569
Rin13_74 in13_73 in13_74 9.241569
Rin13_75 in13_74 in13_75 9.241569
Rin13_76 in13_75 in13_76 9.241569
Rin13_77 in13_76 in13_77 9.241569
Rin13_78 in13_77 in13_78 9.241569
Rin13_79 in13_78 in13_79 9.241569
Rin13_80 in13_79 in13_80 9.241569
Rin13_81 in13_80 in13_81 9.241569
Rin13_82 in13_81 in13_82 9.241569
Rin13_83 in13_82 in13_83 9.241569
Rin13_84 in13_83 in13_84 9.241569
Rin14_1 in14 in14_1 9.241569
Rin14_2 in14_1 in14_2 9.241569
Rin14_3 in14_2 in14_3 9.241569
Rin14_4 in14_3 in14_4 9.241569
Rin14_5 in14_4 in14_5 9.241569
Rin14_6 in14_5 in14_6 9.241569
Rin14_7 in14_6 in14_7 9.241569
Rin14_8 in14_7 in14_8 9.241569
Rin14_9 in14_8 in14_9 9.241569
Rin14_10 in14_9 in14_10 9.241569
Rin14_11 in14_10 in14_11 9.241569
Rin14_12 in14_11 in14_12 9.241569
Rin14_13 in14_12 in14_13 9.241569
Rin14_14 in14_13 in14_14 9.241569
Rin14_15 in14_14 in14_15 9.241569
Rin14_16 in14_15 in14_16 9.241569
Rin14_17 in14_16 in14_17 9.241569
Rin14_18 in14_17 in14_18 9.241569
Rin14_19 in14_18 in14_19 9.241569
Rin14_20 in14_19 in14_20 9.241569
Rin14_21 in14_20 in14_21 9.241569
Rin14_22 in14_21 in14_22 9.241569
Rin14_23 in14_22 in14_23 9.241569
Rin14_24 in14_23 in14_24 9.241569
Rin14_25 in14_24 in14_25 9.241569
Rin14_26 in14_25 in14_26 9.241569
Rin14_27 in14_26 in14_27 9.241569
Rin14_28 in14_27 in14_28 9.241569
Rin14_29 in14 in14_29 9.241569
Rin14_30 in14_29 in14_30 9.241569
Rin14_31 in14_30 in14_31 9.241569
Rin14_32 in14_31 in14_32 9.241569
Rin14_33 in14_32 in14_33 9.241569
Rin14_34 in14_33 in14_34 9.241569
Rin14_35 in14_34 in14_35 9.241569
Rin14_36 in14_35 in14_36 9.241569
Rin14_37 in14_36 in14_37 9.241569
Rin14_38 in14_37 in14_38 9.241569
Rin14_39 in14_38 in14_39 9.241569
Rin14_40 in14_39 in14_40 9.241569
Rin14_41 in14_40 in14_41 9.241569
Rin14_42 in14_41 in14_42 9.241569
Rin14_43 in14_42 in14_43 9.241569
Rin14_44 in14_43 in14_44 9.241569
Rin14_45 in14_44 in14_45 9.241569
Rin14_46 in14_45 in14_46 9.241569
Rin14_47 in14_46 in14_47 9.241569
Rin14_48 in14_47 in14_48 9.241569
Rin14_49 in14_48 in14_49 9.241569
Rin14_50 in14_49 in14_50 9.241569
Rin14_51 in14_50 in14_51 9.241569
Rin14_52 in14_51 in14_52 9.241569
Rin14_53 in14_52 in14_53 9.241569
Rin14_54 in14_53 in14_54 9.241569
Rin14_55 in14_54 in14_55 9.241569
Rin14_56 in14_55 in14_56 9.241569
Rin14_57 in14 in14_57 9.241569
Rin14_58 in14_57 in14_58 9.241569
Rin14_59 in14_58 in14_59 9.241569
Rin14_60 in14_59 in14_60 9.241569
Rin14_61 in14_60 in14_61 9.241569
Rin14_62 in14_61 in14_62 9.241569
Rin14_63 in14_62 in14_63 9.241569
Rin14_64 in14_63 in14_64 9.241569
Rin14_65 in14_64 in14_65 9.241569
Rin14_66 in14_65 in14_66 9.241569
Rin14_67 in14_66 in14_67 9.241569
Rin14_68 in14_67 in14_68 9.241569
Rin14_69 in14_68 in14_69 9.241569
Rin14_70 in14_69 in14_70 9.241569
Rin14_71 in14_70 in14_71 9.241569
Rin14_72 in14_71 in14_72 9.241569
Rin14_73 in14_72 in14_73 9.241569
Rin14_74 in14_73 in14_74 9.241569
Rin14_75 in14_74 in14_75 9.241569
Rin14_76 in14_75 in14_76 9.241569
Rin14_77 in14_76 in14_77 9.241569
Rin14_78 in14_77 in14_78 9.241569
Rin14_79 in14_78 in14_79 9.241569
Rin14_80 in14_79 in14_80 9.241569
Rin14_81 in14_80 in14_81 9.241569
Rin14_82 in14_81 in14_82 9.241569
Rin14_83 in14_82 in14_83 9.241569
Rin14_84 in14_83 in14_84 9.241569
Rin15_1 in15 in15_1 9.241569
Rin15_2 in15_1 in15_2 9.241569
Rin15_3 in15_2 in15_3 9.241569
Rin15_4 in15_3 in15_4 9.241569
Rin15_5 in15_4 in15_5 9.241569
Rin15_6 in15_5 in15_6 9.241569
Rin15_7 in15_6 in15_7 9.241569
Rin15_8 in15_7 in15_8 9.241569
Rin15_9 in15_8 in15_9 9.241569
Rin15_10 in15_9 in15_10 9.241569
Rin15_11 in15_10 in15_11 9.241569
Rin15_12 in15_11 in15_12 9.241569
Rin15_13 in15_12 in15_13 9.241569
Rin15_14 in15_13 in15_14 9.241569
Rin15_15 in15_14 in15_15 9.241569
Rin15_16 in15_15 in15_16 9.241569
Rin15_17 in15_16 in15_17 9.241569
Rin15_18 in15_17 in15_18 9.241569
Rin15_19 in15_18 in15_19 9.241569
Rin15_20 in15_19 in15_20 9.241569
Rin15_21 in15_20 in15_21 9.241569
Rin15_22 in15_21 in15_22 9.241569
Rin15_23 in15_22 in15_23 9.241569
Rin15_24 in15_23 in15_24 9.241569
Rin15_25 in15_24 in15_25 9.241569
Rin15_26 in15_25 in15_26 9.241569
Rin15_27 in15_26 in15_27 9.241569
Rin15_28 in15_27 in15_28 9.241569
Rin15_29 in15 in15_29 9.241569
Rin15_30 in15_29 in15_30 9.241569
Rin15_31 in15_30 in15_31 9.241569
Rin15_32 in15_31 in15_32 9.241569
Rin15_33 in15_32 in15_33 9.241569
Rin15_34 in15_33 in15_34 9.241569
Rin15_35 in15_34 in15_35 9.241569
Rin15_36 in15_35 in15_36 9.241569
Rin15_37 in15_36 in15_37 9.241569
Rin15_38 in15_37 in15_38 9.241569
Rin15_39 in15_38 in15_39 9.241569
Rin15_40 in15_39 in15_40 9.241569
Rin15_41 in15_40 in15_41 9.241569
Rin15_42 in15_41 in15_42 9.241569
Rin15_43 in15_42 in15_43 9.241569
Rin15_44 in15_43 in15_44 9.241569
Rin15_45 in15_44 in15_45 9.241569
Rin15_46 in15_45 in15_46 9.241569
Rin15_47 in15_46 in15_47 9.241569
Rin15_48 in15_47 in15_48 9.241569
Rin15_49 in15_48 in15_49 9.241569
Rin15_50 in15_49 in15_50 9.241569
Rin15_51 in15_50 in15_51 9.241569
Rin15_52 in15_51 in15_52 9.241569
Rin15_53 in15_52 in15_53 9.241569
Rin15_54 in15_53 in15_54 9.241569
Rin15_55 in15_54 in15_55 9.241569
Rin15_56 in15_55 in15_56 9.241569
Rin15_57 in15 in15_57 9.241569
Rin15_58 in15_57 in15_58 9.241569
Rin15_59 in15_58 in15_59 9.241569
Rin15_60 in15_59 in15_60 9.241569
Rin15_61 in15_60 in15_61 9.241569
Rin15_62 in15_61 in15_62 9.241569
Rin15_63 in15_62 in15_63 9.241569
Rin15_64 in15_63 in15_64 9.241569
Rin15_65 in15_64 in15_65 9.241569
Rin15_66 in15_65 in15_66 9.241569
Rin15_67 in15_66 in15_67 9.241569
Rin15_68 in15_67 in15_68 9.241569
Rin15_69 in15_68 in15_69 9.241569
Rin15_70 in15_69 in15_70 9.241569
Rin15_71 in15_70 in15_71 9.241569
Rin15_72 in15_71 in15_72 9.241569
Rin15_73 in15_72 in15_73 9.241569
Rin15_74 in15_73 in15_74 9.241569
Rin15_75 in15_74 in15_75 9.241569
Rin15_76 in15_75 in15_76 9.241569
Rin15_77 in15_76 in15_77 9.241569
Rin15_78 in15_77 in15_78 9.241569
Rin15_79 in15_78 in15_79 9.241569
Rin15_80 in15_79 in15_80 9.241569
Rin15_81 in15_80 in15_81 9.241569
Rin15_82 in15_81 in15_82 9.241569
Rin15_83 in15_82 in15_83 9.241569
Rin15_84 in15_83 in15_84 9.241569
Rin16_1 in16 in16_1 9.241569
Rin16_2 in16_1 in16_2 9.241569
Rin16_3 in16_2 in16_3 9.241569
Rin16_4 in16_3 in16_4 9.241569
Rin16_5 in16_4 in16_5 9.241569
Rin16_6 in16_5 in16_6 9.241569
Rin16_7 in16_6 in16_7 9.241569
Rin16_8 in16_7 in16_8 9.241569
Rin16_9 in16_8 in16_9 9.241569
Rin16_10 in16_9 in16_10 9.241569
Rin16_11 in16_10 in16_11 9.241569
Rin16_12 in16_11 in16_12 9.241569
Rin16_13 in16_12 in16_13 9.241569
Rin16_14 in16_13 in16_14 9.241569
Rin16_15 in16_14 in16_15 9.241569
Rin16_16 in16_15 in16_16 9.241569
Rin16_17 in16_16 in16_17 9.241569
Rin16_18 in16_17 in16_18 9.241569
Rin16_19 in16_18 in16_19 9.241569
Rin16_20 in16_19 in16_20 9.241569
Rin16_21 in16_20 in16_21 9.241569
Rin16_22 in16_21 in16_22 9.241569
Rin16_23 in16_22 in16_23 9.241569
Rin16_24 in16_23 in16_24 9.241569
Rin16_25 in16_24 in16_25 9.241569
Rin16_26 in16_25 in16_26 9.241569
Rin16_27 in16_26 in16_27 9.241569
Rin16_28 in16_27 in16_28 9.241569
Rin16_29 in16 in16_29 9.241569
Rin16_30 in16_29 in16_30 9.241569
Rin16_31 in16_30 in16_31 9.241569
Rin16_32 in16_31 in16_32 9.241569
Rin16_33 in16_32 in16_33 9.241569
Rin16_34 in16_33 in16_34 9.241569
Rin16_35 in16_34 in16_35 9.241569
Rin16_36 in16_35 in16_36 9.241569
Rin16_37 in16_36 in16_37 9.241569
Rin16_38 in16_37 in16_38 9.241569
Rin16_39 in16_38 in16_39 9.241569
Rin16_40 in16_39 in16_40 9.241569
Rin16_41 in16_40 in16_41 9.241569
Rin16_42 in16_41 in16_42 9.241569
Rin16_43 in16_42 in16_43 9.241569
Rin16_44 in16_43 in16_44 9.241569
Rin16_45 in16_44 in16_45 9.241569
Rin16_46 in16_45 in16_46 9.241569
Rin16_47 in16_46 in16_47 9.241569
Rin16_48 in16_47 in16_48 9.241569
Rin16_49 in16_48 in16_49 9.241569
Rin16_50 in16_49 in16_50 9.241569
Rin16_51 in16_50 in16_51 9.241569
Rin16_52 in16_51 in16_52 9.241569
Rin16_53 in16_52 in16_53 9.241569
Rin16_54 in16_53 in16_54 9.241569
Rin16_55 in16_54 in16_55 9.241569
Rin16_56 in16_55 in16_56 9.241569
Rin16_57 in16 in16_57 9.241569
Rin16_58 in16_57 in16_58 9.241569
Rin16_59 in16_58 in16_59 9.241569
Rin16_60 in16_59 in16_60 9.241569
Rin16_61 in16_60 in16_61 9.241569
Rin16_62 in16_61 in16_62 9.241569
Rin16_63 in16_62 in16_63 9.241569
Rin16_64 in16_63 in16_64 9.241569
Rin16_65 in16_64 in16_65 9.241569
Rin16_66 in16_65 in16_66 9.241569
Rin16_67 in16_66 in16_67 9.241569
Rin16_68 in16_67 in16_68 9.241569
Rin16_69 in16_68 in16_69 9.241569
Rin16_70 in16_69 in16_70 9.241569
Rin16_71 in16_70 in16_71 9.241569
Rin16_72 in16_71 in16_72 9.241569
Rin16_73 in16_72 in16_73 9.241569
Rin16_74 in16_73 in16_74 9.241569
Rin16_75 in16_74 in16_75 9.241569
Rin16_76 in16_75 in16_76 9.241569
Rin16_77 in16_76 in16_77 9.241569
Rin16_78 in16_77 in16_78 9.241569
Rin16_79 in16_78 in16_79 9.241569
Rin16_80 in16_79 in16_80 9.241569
Rin16_81 in16_80 in16_81 9.241569
Rin16_82 in16_81 in16_82 9.241569
Rin16_83 in16_82 in16_83 9.241569
Rin16_84 in16_83 in16_84 9.241569
Rin17_1 in17 in17_1 9.241569
Rin17_2 in17_1 in17_2 9.241569
Rin17_3 in17_2 in17_3 9.241569
Rin17_4 in17_3 in17_4 9.241569
Rin17_5 in17_4 in17_5 9.241569
Rin17_6 in17_5 in17_6 9.241569
Rin17_7 in17_6 in17_7 9.241569
Rin17_8 in17_7 in17_8 9.241569
Rin17_9 in17_8 in17_9 9.241569
Rin17_10 in17_9 in17_10 9.241569
Rin17_11 in17_10 in17_11 9.241569
Rin17_12 in17_11 in17_12 9.241569
Rin17_13 in17_12 in17_13 9.241569
Rin17_14 in17_13 in17_14 9.241569
Rin17_15 in17_14 in17_15 9.241569
Rin17_16 in17_15 in17_16 9.241569
Rin17_17 in17_16 in17_17 9.241569
Rin17_18 in17_17 in17_18 9.241569
Rin17_19 in17_18 in17_19 9.241569
Rin17_20 in17_19 in17_20 9.241569
Rin17_21 in17_20 in17_21 9.241569
Rin17_22 in17_21 in17_22 9.241569
Rin17_23 in17_22 in17_23 9.241569
Rin17_24 in17_23 in17_24 9.241569
Rin17_25 in17_24 in17_25 9.241569
Rin17_26 in17_25 in17_26 9.241569
Rin17_27 in17_26 in17_27 9.241569
Rin17_28 in17_27 in17_28 9.241569
Rin17_29 in17 in17_29 9.241569
Rin17_30 in17_29 in17_30 9.241569
Rin17_31 in17_30 in17_31 9.241569
Rin17_32 in17_31 in17_32 9.241569
Rin17_33 in17_32 in17_33 9.241569
Rin17_34 in17_33 in17_34 9.241569
Rin17_35 in17_34 in17_35 9.241569
Rin17_36 in17_35 in17_36 9.241569
Rin17_37 in17_36 in17_37 9.241569
Rin17_38 in17_37 in17_38 9.241569
Rin17_39 in17_38 in17_39 9.241569
Rin17_40 in17_39 in17_40 9.241569
Rin17_41 in17_40 in17_41 9.241569
Rin17_42 in17_41 in17_42 9.241569
Rin17_43 in17_42 in17_43 9.241569
Rin17_44 in17_43 in17_44 9.241569
Rin17_45 in17_44 in17_45 9.241569
Rin17_46 in17_45 in17_46 9.241569
Rin17_47 in17_46 in17_47 9.241569
Rin17_48 in17_47 in17_48 9.241569
Rin17_49 in17_48 in17_49 9.241569
Rin17_50 in17_49 in17_50 9.241569
Rin17_51 in17_50 in17_51 9.241569
Rin17_52 in17_51 in17_52 9.241569
Rin17_53 in17_52 in17_53 9.241569
Rin17_54 in17_53 in17_54 9.241569
Rin17_55 in17_54 in17_55 9.241569
Rin17_56 in17_55 in17_56 9.241569
Rin17_57 in17 in17_57 9.241569
Rin17_58 in17_57 in17_58 9.241569
Rin17_59 in17_58 in17_59 9.241569
Rin17_60 in17_59 in17_60 9.241569
Rin17_61 in17_60 in17_61 9.241569
Rin17_62 in17_61 in17_62 9.241569
Rin17_63 in17_62 in17_63 9.241569
Rin17_64 in17_63 in17_64 9.241569
Rin17_65 in17_64 in17_65 9.241569
Rin17_66 in17_65 in17_66 9.241569
Rin17_67 in17_66 in17_67 9.241569
Rin17_68 in17_67 in17_68 9.241569
Rin17_69 in17_68 in17_69 9.241569
Rin17_70 in17_69 in17_70 9.241569
Rin17_71 in17_70 in17_71 9.241569
Rin17_72 in17_71 in17_72 9.241569
Rin17_73 in17_72 in17_73 9.241569
Rin17_74 in17_73 in17_74 9.241569
Rin17_75 in17_74 in17_75 9.241569
Rin17_76 in17_75 in17_76 9.241569
Rin17_77 in17_76 in17_77 9.241569
Rin17_78 in17_77 in17_78 9.241569
Rin17_79 in17_78 in17_79 9.241569
Rin17_80 in17_79 in17_80 9.241569
Rin17_81 in17_80 in17_81 9.241569
Rin17_82 in17_81 in17_82 9.241569
Rin17_83 in17_82 in17_83 9.241569
Rin17_84 in17_83 in17_84 9.241569
Rin18_1 in18 in18_1 9.241569
Rin18_2 in18_1 in18_2 9.241569
Rin18_3 in18_2 in18_3 9.241569
Rin18_4 in18_3 in18_4 9.241569
Rin18_5 in18_4 in18_5 9.241569
Rin18_6 in18_5 in18_6 9.241569
Rin18_7 in18_6 in18_7 9.241569
Rin18_8 in18_7 in18_8 9.241569
Rin18_9 in18_8 in18_9 9.241569
Rin18_10 in18_9 in18_10 9.241569
Rin18_11 in18_10 in18_11 9.241569
Rin18_12 in18_11 in18_12 9.241569
Rin18_13 in18_12 in18_13 9.241569
Rin18_14 in18_13 in18_14 9.241569
Rin18_15 in18_14 in18_15 9.241569
Rin18_16 in18_15 in18_16 9.241569
Rin18_17 in18_16 in18_17 9.241569
Rin18_18 in18_17 in18_18 9.241569
Rin18_19 in18_18 in18_19 9.241569
Rin18_20 in18_19 in18_20 9.241569
Rin18_21 in18_20 in18_21 9.241569
Rin18_22 in18_21 in18_22 9.241569
Rin18_23 in18_22 in18_23 9.241569
Rin18_24 in18_23 in18_24 9.241569
Rin18_25 in18_24 in18_25 9.241569
Rin18_26 in18_25 in18_26 9.241569
Rin18_27 in18_26 in18_27 9.241569
Rin18_28 in18_27 in18_28 9.241569
Rin18_29 in18 in18_29 9.241569
Rin18_30 in18_29 in18_30 9.241569
Rin18_31 in18_30 in18_31 9.241569
Rin18_32 in18_31 in18_32 9.241569
Rin18_33 in18_32 in18_33 9.241569
Rin18_34 in18_33 in18_34 9.241569
Rin18_35 in18_34 in18_35 9.241569
Rin18_36 in18_35 in18_36 9.241569
Rin18_37 in18_36 in18_37 9.241569
Rin18_38 in18_37 in18_38 9.241569
Rin18_39 in18_38 in18_39 9.241569
Rin18_40 in18_39 in18_40 9.241569
Rin18_41 in18_40 in18_41 9.241569
Rin18_42 in18_41 in18_42 9.241569
Rin18_43 in18_42 in18_43 9.241569
Rin18_44 in18_43 in18_44 9.241569
Rin18_45 in18_44 in18_45 9.241569
Rin18_46 in18_45 in18_46 9.241569
Rin18_47 in18_46 in18_47 9.241569
Rin18_48 in18_47 in18_48 9.241569
Rin18_49 in18_48 in18_49 9.241569
Rin18_50 in18_49 in18_50 9.241569
Rin18_51 in18_50 in18_51 9.241569
Rin18_52 in18_51 in18_52 9.241569
Rin18_53 in18_52 in18_53 9.241569
Rin18_54 in18_53 in18_54 9.241569
Rin18_55 in18_54 in18_55 9.241569
Rin18_56 in18_55 in18_56 9.241569
Rin18_57 in18 in18_57 9.241569
Rin18_58 in18_57 in18_58 9.241569
Rin18_59 in18_58 in18_59 9.241569
Rin18_60 in18_59 in18_60 9.241569
Rin18_61 in18_60 in18_61 9.241569
Rin18_62 in18_61 in18_62 9.241569
Rin18_63 in18_62 in18_63 9.241569
Rin18_64 in18_63 in18_64 9.241569
Rin18_65 in18_64 in18_65 9.241569
Rin18_66 in18_65 in18_66 9.241569
Rin18_67 in18_66 in18_67 9.241569
Rin18_68 in18_67 in18_68 9.241569
Rin18_69 in18_68 in18_69 9.241569
Rin18_70 in18_69 in18_70 9.241569
Rin18_71 in18_70 in18_71 9.241569
Rin18_72 in18_71 in18_72 9.241569
Rin18_73 in18_72 in18_73 9.241569
Rin18_74 in18_73 in18_74 9.241569
Rin18_75 in18_74 in18_75 9.241569
Rin18_76 in18_75 in18_76 9.241569
Rin18_77 in18_76 in18_77 9.241569
Rin18_78 in18_77 in18_78 9.241569
Rin18_79 in18_78 in18_79 9.241569
Rin18_80 in18_79 in18_80 9.241569
Rin18_81 in18_80 in18_81 9.241569
Rin18_82 in18_81 in18_82 9.241569
Rin18_83 in18_82 in18_83 9.241569
Rin18_84 in18_83 in18_84 9.241569
Rin19_1 in19 in19_1 9.241569
Rin19_2 in19_1 in19_2 9.241569
Rin19_3 in19_2 in19_3 9.241569
Rin19_4 in19_3 in19_4 9.241569
Rin19_5 in19_4 in19_5 9.241569
Rin19_6 in19_5 in19_6 9.241569
Rin19_7 in19_6 in19_7 9.241569
Rin19_8 in19_7 in19_8 9.241569
Rin19_9 in19_8 in19_9 9.241569
Rin19_10 in19_9 in19_10 9.241569
Rin19_11 in19_10 in19_11 9.241569
Rin19_12 in19_11 in19_12 9.241569
Rin19_13 in19_12 in19_13 9.241569
Rin19_14 in19_13 in19_14 9.241569
Rin19_15 in19_14 in19_15 9.241569
Rin19_16 in19_15 in19_16 9.241569
Rin19_17 in19_16 in19_17 9.241569
Rin19_18 in19_17 in19_18 9.241569
Rin19_19 in19_18 in19_19 9.241569
Rin19_20 in19_19 in19_20 9.241569
Rin19_21 in19_20 in19_21 9.241569
Rin19_22 in19_21 in19_22 9.241569
Rin19_23 in19_22 in19_23 9.241569
Rin19_24 in19_23 in19_24 9.241569
Rin19_25 in19_24 in19_25 9.241569
Rin19_26 in19_25 in19_26 9.241569
Rin19_27 in19_26 in19_27 9.241569
Rin19_28 in19_27 in19_28 9.241569
Rin19_29 in19 in19_29 9.241569
Rin19_30 in19_29 in19_30 9.241569
Rin19_31 in19_30 in19_31 9.241569
Rin19_32 in19_31 in19_32 9.241569
Rin19_33 in19_32 in19_33 9.241569
Rin19_34 in19_33 in19_34 9.241569
Rin19_35 in19_34 in19_35 9.241569
Rin19_36 in19_35 in19_36 9.241569
Rin19_37 in19_36 in19_37 9.241569
Rin19_38 in19_37 in19_38 9.241569
Rin19_39 in19_38 in19_39 9.241569
Rin19_40 in19_39 in19_40 9.241569
Rin19_41 in19_40 in19_41 9.241569
Rin19_42 in19_41 in19_42 9.241569
Rin19_43 in19_42 in19_43 9.241569
Rin19_44 in19_43 in19_44 9.241569
Rin19_45 in19_44 in19_45 9.241569
Rin19_46 in19_45 in19_46 9.241569
Rin19_47 in19_46 in19_47 9.241569
Rin19_48 in19_47 in19_48 9.241569
Rin19_49 in19_48 in19_49 9.241569
Rin19_50 in19_49 in19_50 9.241569
Rin19_51 in19_50 in19_51 9.241569
Rin19_52 in19_51 in19_52 9.241569
Rin19_53 in19_52 in19_53 9.241569
Rin19_54 in19_53 in19_54 9.241569
Rin19_55 in19_54 in19_55 9.241569
Rin19_56 in19_55 in19_56 9.241569
Rin19_57 in19 in19_57 9.241569
Rin19_58 in19_57 in19_58 9.241569
Rin19_59 in19_58 in19_59 9.241569
Rin19_60 in19_59 in19_60 9.241569
Rin19_61 in19_60 in19_61 9.241569
Rin19_62 in19_61 in19_62 9.241569
Rin19_63 in19_62 in19_63 9.241569
Rin19_64 in19_63 in19_64 9.241569
Rin19_65 in19_64 in19_65 9.241569
Rin19_66 in19_65 in19_66 9.241569
Rin19_67 in19_66 in19_67 9.241569
Rin19_68 in19_67 in19_68 9.241569
Rin19_69 in19_68 in19_69 9.241569
Rin19_70 in19_69 in19_70 9.241569
Rin19_71 in19_70 in19_71 9.241569
Rin19_72 in19_71 in19_72 9.241569
Rin19_73 in19_72 in19_73 9.241569
Rin19_74 in19_73 in19_74 9.241569
Rin19_75 in19_74 in19_75 9.241569
Rin19_76 in19_75 in19_76 9.241569
Rin19_77 in19_76 in19_77 9.241569
Rin19_78 in19_77 in19_78 9.241569
Rin19_79 in19_78 in19_79 9.241569
Rin19_80 in19_79 in19_80 9.241569
Rin19_81 in19_80 in19_81 9.241569
Rin19_82 in19_81 in19_82 9.241569
Rin19_83 in19_82 in19_83 9.241569
Rin19_84 in19_83 in19_84 9.241569
Rin20_1 in20 in20_1 9.241569
Rin20_2 in20_1 in20_2 9.241569
Rin20_3 in20_2 in20_3 9.241569
Rin20_4 in20_3 in20_4 9.241569
Rin20_5 in20_4 in20_5 9.241569
Rin20_6 in20_5 in20_6 9.241569
Rin20_7 in20_6 in20_7 9.241569
Rin20_8 in20_7 in20_8 9.241569
Rin20_9 in20_8 in20_9 9.241569
Rin20_10 in20_9 in20_10 9.241569
Rin20_11 in20_10 in20_11 9.241569
Rin20_12 in20_11 in20_12 9.241569
Rin20_13 in20_12 in20_13 9.241569
Rin20_14 in20_13 in20_14 9.241569
Rin20_15 in20_14 in20_15 9.241569
Rin20_16 in20_15 in20_16 9.241569
Rin20_17 in20_16 in20_17 9.241569
Rin20_18 in20_17 in20_18 9.241569
Rin20_19 in20_18 in20_19 9.241569
Rin20_20 in20_19 in20_20 9.241569
Rin20_21 in20_20 in20_21 9.241569
Rin20_22 in20_21 in20_22 9.241569
Rin20_23 in20_22 in20_23 9.241569
Rin20_24 in20_23 in20_24 9.241569
Rin20_25 in20_24 in20_25 9.241569
Rin20_26 in20_25 in20_26 9.241569
Rin20_27 in20_26 in20_27 9.241569
Rin20_28 in20_27 in20_28 9.241569
Rin20_29 in20 in20_29 9.241569
Rin20_30 in20_29 in20_30 9.241569
Rin20_31 in20_30 in20_31 9.241569
Rin20_32 in20_31 in20_32 9.241569
Rin20_33 in20_32 in20_33 9.241569
Rin20_34 in20_33 in20_34 9.241569
Rin20_35 in20_34 in20_35 9.241569
Rin20_36 in20_35 in20_36 9.241569
Rin20_37 in20_36 in20_37 9.241569
Rin20_38 in20_37 in20_38 9.241569
Rin20_39 in20_38 in20_39 9.241569
Rin20_40 in20_39 in20_40 9.241569
Rin20_41 in20_40 in20_41 9.241569
Rin20_42 in20_41 in20_42 9.241569
Rin20_43 in20_42 in20_43 9.241569
Rin20_44 in20_43 in20_44 9.241569
Rin20_45 in20_44 in20_45 9.241569
Rin20_46 in20_45 in20_46 9.241569
Rin20_47 in20_46 in20_47 9.241569
Rin20_48 in20_47 in20_48 9.241569
Rin20_49 in20_48 in20_49 9.241569
Rin20_50 in20_49 in20_50 9.241569
Rin20_51 in20_50 in20_51 9.241569
Rin20_52 in20_51 in20_52 9.241569
Rin20_53 in20_52 in20_53 9.241569
Rin20_54 in20_53 in20_54 9.241569
Rin20_55 in20_54 in20_55 9.241569
Rin20_56 in20_55 in20_56 9.241569
Rin20_57 in20 in20_57 9.241569
Rin20_58 in20_57 in20_58 9.241569
Rin20_59 in20_58 in20_59 9.241569
Rin20_60 in20_59 in20_60 9.241569
Rin20_61 in20_60 in20_61 9.241569
Rin20_62 in20_61 in20_62 9.241569
Rin20_63 in20_62 in20_63 9.241569
Rin20_64 in20_63 in20_64 9.241569
Rin20_65 in20_64 in20_65 9.241569
Rin20_66 in20_65 in20_66 9.241569
Rin20_67 in20_66 in20_67 9.241569
Rin20_68 in20_67 in20_68 9.241569
Rin20_69 in20_68 in20_69 9.241569
Rin20_70 in20_69 in20_70 9.241569
Rin20_71 in20_70 in20_71 9.241569
Rin20_72 in20_71 in20_72 9.241569
Rin20_73 in20_72 in20_73 9.241569
Rin20_74 in20_73 in20_74 9.241569
Rin20_75 in20_74 in20_75 9.241569
Rin20_76 in20_75 in20_76 9.241569
Rin20_77 in20_76 in20_77 9.241569
Rin20_78 in20_77 in20_78 9.241569
Rin20_79 in20_78 in20_79 9.241569
Rin20_80 in20_79 in20_80 9.241569
Rin20_81 in20_80 in20_81 9.241569
Rin20_82 in20_81 in20_82 9.241569
Rin20_83 in20_82 in20_83 9.241569
Rin20_84 in20_83 in20_84 9.241569
Rin21_1 in21 in21_1 9.241569
Rin21_2 in21_1 in21_2 9.241569
Rin21_3 in21_2 in21_3 9.241569
Rin21_4 in21_3 in21_4 9.241569
Rin21_5 in21_4 in21_5 9.241569
Rin21_6 in21_5 in21_6 9.241569
Rin21_7 in21_6 in21_7 9.241569
Rin21_8 in21_7 in21_8 9.241569
Rin21_9 in21_8 in21_9 9.241569
Rin21_10 in21_9 in21_10 9.241569
Rin21_11 in21_10 in21_11 9.241569
Rin21_12 in21_11 in21_12 9.241569
Rin21_13 in21_12 in21_13 9.241569
Rin21_14 in21_13 in21_14 9.241569
Rin21_15 in21_14 in21_15 9.241569
Rin21_16 in21_15 in21_16 9.241569
Rin21_17 in21_16 in21_17 9.241569
Rin21_18 in21_17 in21_18 9.241569
Rin21_19 in21_18 in21_19 9.241569
Rin21_20 in21_19 in21_20 9.241569
Rin21_21 in21_20 in21_21 9.241569
Rin21_22 in21_21 in21_22 9.241569
Rin21_23 in21_22 in21_23 9.241569
Rin21_24 in21_23 in21_24 9.241569
Rin21_25 in21_24 in21_25 9.241569
Rin21_26 in21_25 in21_26 9.241569
Rin21_27 in21_26 in21_27 9.241569
Rin21_28 in21_27 in21_28 9.241569
Rin21_29 in21 in21_29 9.241569
Rin21_30 in21_29 in21_30 9.241569
Rin21_31 in21_30 in21_31 9.241569
Rin21_32 in21_31 in21_32 9.241569
Rin21_33 in21_32 in21_33 9.241569
Rin21_34 in21_33 in21_34 9.241569
Rin21_35 in21_34 in21_35 9.241569
Rin21_36 in21_35 in21_36 9.241569
Rin21_37 in21_36 in21_37 9.241569
Rin21_38 in21_37 in21_38 9.241569
Rin21_39 in21_38 in21_39 9.241569
Rin21_40 in21_39 in21_40 9.241569
Rin21_41 in21_40 in21_41 9.241569
Rin21_42 in21_41 in21_42 9.241569
Rin21_43 in21_42 in21_43 9.241569
Rin21_44 in21_43 in21_44 9.241569
Rin21_45 in21_44 in21_45 9.241569
Rin21_46 in21_45 in21_46 9.241569
Rin21_47 in21_46 in21_47 9.241569
Rin21_48 in21_47 in21_48 9.241569
Rin21_49 in21_48 in21_49 9.241569
Rin21_50 in21_49 in21_50 9.241569
Rin21_51 in21_50 in21_51 9.241569
Rin21_52 in21_51 in21_52 9.241569
Rin21_53 in21_52 in21_53 9.241569
Rin21_54 in21_53 in21_54 9.241569
Rin21_55 in21_54 in21_55 9.241569
Rin21_56 in21_55 in21_56 9.241569
Rin21_57 in21 in21_57 9.241569
Rin21_58 in21_57 in21_58 9.241569
Rin21_59 in21_58 in21_59 9.241569
Rin21_60 in21_59 in21_60 9.241569
Rin21_61 in21_60 in21_61 9.241569
Rin21_62 in21_61 in21_62 9.241569
Rin21_63 in21_62 in21_63 9.241569
Rin21_64 in21_63 in21_64 9.241569
Rin21_65 in21_64 in21_65 9.241569
Rin21_66 in21_65 in21_66 9.241569
Rin21_67 in21_66 in21_67 9.241569
Rin21_68 in21_67 in21_68 9.241569
Rin21_69 in21_68 in21_69 9.241569
Rin21_70 in21_69 in21_70 9.241569
Rin21_71 in21_70 in21_71 9.241569
Rin21_72 in21_71 in21_72 9.241569
Rin21_73 in21_72 in21_73 9.241569
Rin21_74 in21_73 in21_74 9.241569
Rin21_75 in21_74 in21_75 9.241569
Rin21_76 in21_75 in21_76 9.241569
Rin21_77 in21_76 in21_77 9.241569
Rin21_78 in21_77 in21_78 9.241569
Rin21_79 in21_78 in21_79 9.241569
Rin21_80 in21_79 in21_80 9.241569
Rin21_81 in21_80 in21_81 9.241569
Rin21_82 in21_81 in21_82 9.241569
Rin21_83 in21_82 in21_83 9.241569
Rin21_84 in21_83 in21_84 9.241569
Rin22_1 in22 in22_1 9.241569
Rin22_2 in22_1 in22_2 9.241569
Rin22_3 in22_2 in22_3 9.241569
Rin22_4 in22_3 in22_4 9.241569
Rin22_5 in22_4 in22_5 9.241569
Rin22_6 in22_5 in22_6 9.241569
Rin22_7 in22_6 in22_7 9.241569
Rin22_8 in22_7 in22_8 9.241569
Rin22_9 in22_8 in22_9 9.241569
Rin22_10 in22_9 in22_10 9.241569
Rin22_11 in22_10 in22_11 9.241569
Rin22_12 in22_11 in22_12 9.241569
Rin22_13 in22_12 in22_13 9.241569
Rin22_14 in22_13 in22_14 9.241569
Rin22_15 in22_14 in22_15 9.241569
Rin22_16 in22_15 in22_16 9.241569
Rin22_17 in22_16 in22_17 9.241569
Rin22_18 in22_17 in22_18 9.241569
Rin22_19 in22_18 in22_19 9.241569
Rin22_20 in22_19 in22_20 9.241569
Rin22_21 in22_20 in22_21 9.241569
Rin22_22 in22_21 in22_22 9.241569
Rin22_23 in22_22 in22_23 9.241569
Rin22_24 in22_23 in22_24 9.241569
Rin22_25 in22_24 in22_25 9.241569
Rin22_26 in22_25 in22_26 9.241569
Rin22_27 in22_26 in22_27 9.241569
Rin22_28 in22_27 in22_28 9.241569
Rin22_29 in22 in22_29 9.241569
Rin22_30 in22_29 in22_30 9.241569
Rin22_31 in22_30 in22_31 9.241569
Rin22_32 in22_31 in22_32 9.241569
Rin22_33 in22_32 in22_33 9.241569
Rin22_34 in22_33 in22_34 9.241569
Rin22_35 in22_34 in22_35 9.241569
Rin22_36 in22_35 in22_36 9.241569
Rin22_37 in22_36 in22_37 9.241569
Rin22_38 in22_37 in22_38 9.241569
Rin22_39 in22_38 in22_39 9.241569
Rin22_40 in22_39 in22_40 9.241569
Rin22_41 in22_40 in22_41 9.241569
Rin22_42 in22_41 in22_42 9.241569
Rin22_43 in22_42 in22_43 9.241569
Rin22_44 in22_43 in22_44 9.241569
Rin22_45 in22_44 in22_45 9.241569
Rin22_46 in22_45 in22_46 9.241569
Rin22_47 in22_46 in22_47 9.241569
Rin22_48 in22_47 in22_48 9.241569
Rin22_49 in22_48 in22_49 9.241569
Rin22_50 in22_49 in22_50 9.241569
Rin22_51 in22_50 in22_51 9.241569
Rin22_52 in22_51 in22_52 9.241569
Rin22_53 in22_52 in22_53 9.241569
Rin22_54 in22_53 in22_54 9.241569
Rin22_55 in22_54 in22_55 9.241569
Rin22_56 in22_55 in22_56 9.241569
Rin22_57 in22 in22_57 9.241569
Rin22_58 in22_57 in22_58 9.241569
Rin22_59 in22_58 in22_59 9.241569
Rin22_60 in22_59 in22_60 9.241569
Rin22_61 in22_60 in22_61 9.241569
Rin22_62 in22_61 in22_62 9.241569
Rin22_63 in22_62 in22_63 9.241569
Rin22_64 in22_63 in22_64 9.241569
Rin22_65 in22_64 in22_65 9.241569
Rin22_66 in22_65 in22_66 9.241569
Rin22_67 in22_66 in22_67 9.241569
Rin22_68 in22_67 in22_68 9.241569
Rin22_69 in22_68 in22_69 9.241569
Rin22_70 in22_69 in22_70 9.241569
Rin22_71 in22_70 in22_71 9.241569
Rin22_72 in22_71 in22_72 9.241569
Rin22_73 in22_72 in22_73 9.241569
Rin22_74 in22_73 in22_74 9.241569
Rin22_75 in22_74 in22_75 9.241569
Rin22_76 in22_75 in22_76 9.241569
Rin22_77 in22_76 in22_77 9.241569
Rin22_78 in22_77 in22_78 9.241569
Rin22_79 in22_78 in22_79 9.241569
Rin22_80 in22_79 in22_80 9.241569
Rin22_81 in22_80 in22_81 9.241569
Rin22_82 in22_81 in22_82 9.241569
Rin22_83 in22_82 in22_83 9.241569
Rin22_84 in22_83 in22_84 9.241569
Rin23_1 in23 in23_1 9.241569
Rin23_2 in23_1 in23_2 9.241569
Rin23_3 in23_2 in23_3 9.241569
Rin23_4 in23_3 in23_4 9.241569
Rin23_5 in23_4 in23_5 9.241569
Rin23_6 in23_5 in23_6 9.241569
Rin23_7 in23_6 in23_7 9.241569
Rin23_8 in23_7 in23_8 9.241569
Rin23_9 in23_8 in23_9 9.241569
Rin23_10 in23_9 in23_10 9.241569
Rin23_11 in23_10 in23_11 9.241569
Rin23_12 in23_11 in23_12 9.241569
Rin23_13 in23_12 in23_13 9.241569
Rin23_14 in23_13 in23_14 9.241569
Rin23_15 in23_14 in23_15 9.241569
Rin23_16 in23_15 in23_16 9.241569
Rin23_17 in23_16 in23_17 9.241569
Rin23_18 in23_17 in23_18 9.241569
Rin23_19 in23_18 in23_19 9.241569
Rin23_20 in23_19 in23_20 9.241569
Rin23_21 in23_20 in23_21 9.241569
Rin23_22 in23_21 in23_22 9.241569
Rin23_23 in23_22 in23_23 9.241569
Rin23_24 in23_23 in23_24 9.241569
Rin23_25 in23_24 in23_25 9.241569
Rin23_26 in23_25 in23_26 9.241569
Rin23_27 in23_26 in23_27 9.241569
Rin23_28 in23_27 in23_28 9.241569
Rin23_29 in23 in23_29 9.241569
Rin23_30 in23_29 in23_30 9.241569
Rin23_31 in23_30 in23_31 9.241569
Rin23_32 in23_31 in23_32 9.241569
Rin23_33 in23_32 in23_33 9.241569
Rin23_34 in23_33 in23_34 9.241569
Rin23_35 in23_34 in23_35 9.241569
Rin23_36 in23_35 in23_36 9.241569
Rin23_37 in23_36 in23_37 9.241569
Rin23_38 in23_37 in23_38 9.241569
Rin23_39 in23_38 in23_39 9.241569
Rin23_40 in23_39 in23_40 9.241569
Rin23_41 in23_40 in23_41 9.241569
Rin23_42 in23_41 in23_42 9.241569
Rin23_43 in23_42 in23_43 9.241569
Rin23_44 in23_43 in23_44 9.241569
Rin23_45 in23_44 in23_45 9.241569
Rin23_46 in23_45 in23_46 9.241569
Rin23_47 in23_46 in23_47 9.241569
Rin23_48 in23_47 in23_48 9.241569
Rin23_49 in23_48 in23_49 9.241569
Rin23_50 in23_49 in23_50 9.241569
Rin23_51 in23_50 in23_51 9.241569
Rin23_52 in23_51 in23_52 9.241569
Rin23_53 in23_52 in23_53 9.241569
Rin23_54 in23_53 in23_54 9.241569
Rin23_55 in23_54 in23_55 9.241569
Rin23_56 in23_55 in23_56 9.241569
Rin23_57 in23 in23_57 9.241569
Rin23_58 in23_57 in23_58 9.241569
Rin23_59 in23_58 in23_59 9.241569
Rin23_60 in23_59 in23_60 9.241569
Rin23_61 in23_60 in23_61 9.241569
Rin23_62 in23_61 in23_62 9.241569
Rin23_63 in23_62 in23_63 9.241569
Rin23_64 in23_63 in23_64 9.241569
Rin23_65 in23_64 in23_65 9.241569
Rin23_66 in23_65 in23_66 9.241569
Rin23_67 in23_66 in23_67 9.241569
Rin23_68 in23_67 in23_68 9.241569
Rin23_69 in23_68 in23_69 9.241569
Rin23_70 in23_69 in23_70 9.241569
Rin23_71 in23_70 in23_71 9.241569
Rin23_72 in23_71 in23_72 9.241569
Rin23_73 in23_72 in23_73 9.241569
Rin23_74 in23_73 in23_74 9.241569
Rin23_75 in23_74 in23_75 9.241569
Rin23_76 in23_75 in23_76 9.241569
Rin23_77 in23_76 in23_77 9.241569
Rin23_78 in23_77 in23_78 9.241569
Rin23_79 in23_78 in23_79 9.241569
Rin23_80 in23_79 in23_80 9.241569
Rin23_81 in23_80 in23_81 9.241569
Rin23_82 in23_81 in23_82 9.241569
Rin23_83 in23_82 in23_83 9.241569
Rin23_84 in23_83 in23_84 9.241569
Rin24_1 in24 in24_1 9.241569
Rin24_2 in24_1 in24_2 9.241569
Rin24_3 in24_2 in24_3 9.241569
Rin24_4 in24_3 in24_4 9.241569
Rin24_5 in24_4 in24_5 9.241569
Rin24_6 in24_5 in24_6 9.241569
Rin24_7 in24_6 in24_7 9.241569
Rin24_8 in24_7 in24_8 9.241569
Rin24_9 in24_8 in24_9 9.241569
Rin24_10 in24_9 in24_10 9.241569
Rin24_11 in24_10 in24_11 9.241569
Rin24_12 in24_11 in24_12 9.241569
Rin24_13 in24_12 in24_13 9.241569
Rin24_14 in24_13 in24_14 9.241569
Rin24_15 in24_14 in24_15 9.241569
Rin24_16 in24_15 in24_16 9.241569
Rin24_17 in24_16 in24_17 9.241569
Rin24_18 in24_17 in24_18 9.241569
Rin24_19 in24_18 in24_19 9.241569
Rin24_20 in24_19 in24_20 9.241569
Rin24_21 in24_20 in24_21 9.241569
Rin24_22 in24_21 in24_22 9.241569
Rin24_23 in24_22 in24_23 9.241569
Rin24_24 in24_23 in24_24 9.241569
Rin24_25 in24_24 in24_25 9.241569
Rin24_26 in24_25 in24_26 9.241569
Rin24_27 in24_26 in24_27 9.241569
Rin24_28 in24_27 in24_28 9.241569
Rin24_29 in24 in24_29 9.241569
Rin24_30 in24_29 in24_30 9.241569
Rin24_31 in24_30 in24_31 9.241569
Rin24_32 in24_31 in24_32 9.241569
Rin24_33 in24_32 in24_33 9.241569
Rin24_34 in24_33 in24_34 9.241569
Rin24_35 in24_34 in24_35 9.241569
Rin24_36 in24_35 in24_36 9.241569
Rin24_37 in24_36 in24_37 9.241569
Rin24_38 in24_37 in24_38 9.241569
Rin24_39 in24_38 in24_39 9.241569
Rin24_40 in24_39 in24_40 9.241569
Rin24_41 in24_40 in24_41 9.241569
Rin24_42 in24_41 in24_42 9.241569
Rin24_43 in24_42 in24_43 9.241569
Rin24_44 in24_43 in24_44 9.241569
Rin24_45 in24_44 in24_45 9.241569
Rin24_46 in24_45 in24_46 9.241569
Rin24_47 in24_46 in24_47 9.241569
Rin24_48 in24_47 in24_48 9.241569
Rin24_49 in24_48 in24_49 9.241569
Rin24_50 in24_49 in24_50 9.241569
Rin24_51 in24_50 in24_51 9.241569
Rin24_52 in24_51 in24_52 9.241569
Rin24_53 in24_52 in24_53 9.241569
Rin24_54 in24_53 in24_54 9.241569
Rin24_55 in24_54 in24_55 9.241569
Rin24_56 in24_55 in24_56 9.241569
Rin24_57 in24 in24_57 9.241569
Rin24_58 in24_57 in24_58 9.241569
Rin24_59 in24_58 in24_59 9.241569
Rin24_60 in24_59 in24_60 9.241569
Rin24_61 in24_60 in24_61 9.241569
Rin24_62 in24_61 in24_62 9.241569
Rin24_63 in24_62 in24_63 9.241569
Rin24_64 in24_63 in24_64 9.241569
Rin24_65 in24_64 in24_65 9.241569
Rin24_66 in24_65 in24_66 9.241569
Rin24_67 in24_66 in24_67 9.241569
Rin24_68 in24_67 in24_68 9.241569
Rin24_69 in24_68 in24_69 9.241569
Rin24_70 in24_69 in24_70 9.241569
Rin24_71 in24_70 in24_71 9.241569
Rin24_72 in24_71 in24_72 9.241569
Rin24_73 in24_72 in24_73 9.241569
Rin24_74 in24_73 in24_74 9.241569
Rin24_75 in24_74 in24_75 9.241569
Rin24_76 in24_75 in24_76 9.241569
Rin24_77 in24_76 in24_77 9.241569
Rin24_78 in24_77 in24_78 9.241569
Rin24_79 in24_78 in24_79 9.241569
Rin24_80 in24_79 in24_80 9.241569
Rin24_81 in24_80 in24_81 9.241569
Rin24_82 in24_81 in24_82 9.241569
Rin24_83 in24_82 in24_83 9.241569
Rin24_84 in24_83 in24_84 9.241569
Rin25_1 in25 in25_1 9.241569
Rin25_2 in25_1 in25_2 9.241569
Rin25_3 in25_2 in25_3 9.241569
Rin25_4 in25_3 in25_4 9.241569
Rin25_5 in25_4 in25_5 9.241569
Rin25_6 in25_5 in25_6 9.241569
Rin25_7 in25_6 in25_7 9.241569
Rin25_8 in25_7 in25_8 9.241569
Rin25_9 in25_8 in25_9 9.241569
Rin25_10 in25_9 in25_10 9.241569
Rin25_11 in25_10 in25_11 9.241569
Rin25_12 in25_11 in25_12 9.241569
Rin25_13 in25_12 in25_13 9.241569
Rin25_14 in25_13 in25_14 9.241569
Rin25_15 in25_14 in25_15 9.241569
Rin25_16 in25_15 in25_16 9.241569
Rin25_17 in25_16 in25_17 9.241569
Rin25_18 in25_17 in25_18 9.241569
Rin25_19 in25_18 in25_19 9.241569
Rin25_20 in25_19 in25_20 9.241569
Rin25_21 in25_20 in25_21 9.241569
Rin25_22 in25_21 in25_22 9.241569
Rin25_23 in25_22 in25_23 9.241569
Rin25_24 in25_23 in25_24 9.241569
Rin25_25 in25_24 in25_25 9.241569
Rin25_26 in25_25 in25_26 9.241569
Rin25_27 in25_26 in25_27 9.241569
Rin25_28 in25_27 in25_28 9.241569
Rin25_29 in25 in25_29 9.241569
Rin25_30 in25_29 in25_30 9.241569
Rin25_31 in25_30 in25_31 9.241569
Rin25_32 in25_31 in25_32 9.241569
Rin25_33 in25_32 in25_33 9.241569
Rin25_34 in25_33 in25_34 9.241569
Rin25_35 in25_34 in25_35 9.241569
Rin25_36 in25_35 in25_36 9.241569
Rin25_37 in25_36 in25_37 9.241569
Rin25_38 in25_37 in25_38 9.241569
Rin25_39 in25_38 in25_39 9.241569
Rin25_40 in25_39 in25_40 9.241569
Rin25_41 in25_40 in25_41 9.241569
Rin25_42 in25_41 in25_42 9.241569
Rin25_43 in25_42 in25_43 9.241569
Rin25_44 in25_43 in25_44 9.241569
Rin25_45 in25_44 in25_45 9.241569
Rin25_46 in25_45 in25_46 9.241569
Rin25_47 in25_46 in25_47 9.241569
Rin25_48 in25_47 in25_48 9.241569
Rin25_49 in25_48 in25_49 9.241569
Rin25_50 in25_49 in25_50 9.241569
Rin25_51 in25_50 in25_51 9.241569
Rin25_52 in25_51 in25_52 9.241569
Rin25_53 in25_52 in25_53 9.241569
Rin25_54 in25_53 in25_54 9.241569
Rin25_55 in25_54 in25_55 9.241569
Rin25_56 in25_55 in25_56 9.241569
Rin25_57 in25 in25_57 9.241569
Rin25_58 in25_57 in25_58 9.241569
Rin25_59 in25_58 in25_59 9.241569
Rin25_60 in25_59 in25_60 9.241569
Rin25_61 in25_60 in25_61 9.241569
Rin25_62 in25_61 in25_62 9.241569
Rin25_63 in25_62 in25_63 9.241569
Rin25_64 in25_63 in25_64 9.241569
Rin25_65 in25_64 in25_65 9.241569
Rin25_66 in25_65 in25_66 9.241569
Rin25_67 in25_66 in25_67 9.241569
Rin25_68 in25_67 in25_68 9.241569
Rin25_69 in25_68 in25_69 9.241569
Rin25_70 in25_69 in25_70 9.241569
Rin25_71 in25_70 in25_71 9.241569
Rin25_72 in25_71 in25_72 9.241569
Rin25_73 in25_72 in25_73 9.241569
Rin25_74 in25_73 in25_74 9.241569
Rin25_75 in25_74 in25_75 9.241569
Rin25_76 in25_75 in25_76 9.241569
Rin25_77 in25_76 in25_77 9.241569
Rin25_78 in25_77 in25_78 9.241569
Rin25_79 in25_78 in25_79 9.241569
Rin25_80 in25_79 in25_80 9.241569
Rin25_81 in25_80 in25_81 9.241569
Rin25_82 in25_81 in25_82 9.241569
Rin25_83 in25_82 in25_83 9.241569
Rin25_84 in25_83 in25_84 9.241569
Rin26_1 in26 in26_1 9.241569
Rin26_2 in26_1 in26_2 9.241569
Rin26_3 in26_2 in26_3 9.241569
Rin26_4 in26_3 in26_4 9.241569
Rin26_5 in26_4 in26_5 9.241569
Rin26_6 in26_5 in26_6 9.241569
Rin26_7 in26_6 in26_7 9.241569
Rin26_8 in26_7 in26_8 9.241569
Rin26_9 in26_8 in26_9 9.241569
Rin26_10 in26_9 in26_10 9.241569
Rin26_11 in26_10 in26_11 9.241569
Rin26_12 in26_11 in26_12 9.241569
Rin26_13 in26_12 in26_13 9.241569
Rin26_14 in26_13 in26_14 9.241569
Rin26_15 in26_14 in26_15 9.241569
Rin26_16 in26_15 in26_16 9.241569
Rin26_17 in26_16 in26_17 9.241569
Rin26_18 in26_17 in26_18 9.241569
Rin26_19 in26_18 in26_19 9.241569
Rin26_20 in26_19 in26_20 9.241569
Rin26_21 in26_20 in26_21 9.241569
Rin26_22 in26_21 in26_22 9.241569
Rin26_23 in26_22 in26_23 9.241569
Rin26_24 in26_23 in26_24 9.241569
Rin26_25 in26_24 in26_25 9.241569
Rin26_26 in26_25 in26_26 9.241569
Rin26_27 in26_26 in26_27 9.241569
Rin26_28 in26_27 in26_28 9.241569
Rin26_29 in26 in26_29 9.241569
Rin26_30 in26_29 in26_30 9.241569
Rin26_31 in26_30 in26_31 9.241569
Rin26_32 in26_31 in26_32 9.241569
Rin26_33 in26_32 in26_33 9.241569
Rin26_34 in26_33 in26_34 9.241569
Rin26_35 in26_34 in26_35 9.241569
Rin26_36 in26_35 in26_36 9.241569
Rin26_37 in26_36 in26_37 9.241569
Rin26_38 in26_37 in26_38 9.241569
Rin26_39 in26_38 in26_39 9.241569
Rin26_40 in26_39 in26_40 9.241569
Rin26_41 in26_40 in26_41 9.241569
Rin26_42 in26_41 in26_42 9.241569
Rin26_43 in26_42 in26_43 9.241569
Rin26_44 in26_43 in26_44 9.241569
Rin26_45 in26_44 in26_45 9.241569
Rin26_46 in26_45 in26_46 9.241569
Rin26_47 in26_46 in26_47 9.241569
Rin26_48 in26_47 in26_48 9.241569
Rin26_49 in26_48 in26_49 9.241569
Rin26_50 in26_49 in26_50 9.241569
Rin26_51 in26_50 in26_51 9.241569
Rin26_52 in26_51 in26_52 9.241569
Rin26_53 in26_52 in26_53 9.241569
Rin26_54 in26_53 in26_54 9.241569
Rin26_55 in26_54 in26_55 9.241569
Rin26_56 in26_55 in26_56 9.241569
Rin26_57 in26 in26_57 9.241569
Rin26_58 in26_57 in26_58 9.241569
Rin26_59 in26_58 in26_59 9.241569
Rin26_60 in26_59 in26_60 9.241569
Rin26_61 in26_60 in26_61 9.241569
Rin26_62 in26_61 in26_62 9.241569
Rin26_63 in26_62 in26_63 9.241569
Rin26_64 in26_63 in26_64 9.241569
Rin26_65 in26_64 in26_65 9.241569
Rin26_66 in26_65 in26_66 9.241569
Rin26_67 in26_66 in26_67 9.241569
Rin26_68 in26_67 in26_68 9.241569
Rin26_69 in26_68 in26_69 9.241569
Rin26_70 in26_69 in26_70 9.241569
Rin26_71 in26_70 in26_71 9.241569
Rin26_72 in26_71 in26_72 9.241569
Rin26_73 in26_72 in26_73 9.241569
Rin26_74 in26_73 in26_74 9.241569
Rin26_75 in26_74 in26_75 9.241569
Rin26_76 in26_75 in26_76 9.241569
Rin26_77 in26_76 in26_77 9.241569
Rin26_78 in26_77 in26_78 9.241569
Rin26_79 in26_78 in26_79 9.241569
Rin26_80 in26_79 in26_80 9.241569
Rin26_81 in26_80 in26_81 9.241569
Rin26_82 in26_81 in26_82 9.241569
Rin26_83 in26_82 in26_83 9.241569
Rin26_84 in26_83 in26_84 9.241569
Rin27_1 in27 in27_1 9.241569
Rin27_2 in27_1 in27_2 9.241569
Rin27_3 in27_2 in27_3 9.241569
Rin27_4 in27_3 in27_4 9.241569
Rin27_5 in27_4 in27_5 9.241569
Rin27_6 in27_5 in27_6 9.241569
Rin27_7 in27_6 in27_7 9.241569
Rin27_8 in27_7 in27_8 9.241569
Rin27_9 in27_8 in27_9 9.241569
Rin27_10 in27_9 in27_10 9.241569
Rin27_11 in27_10 in27_11 9.241569
Rin27_12 in27_11 in27_12 9.241569
Rin27_13 in27_12 in27_13 9.241569
Rin27_14 in27_13 in27_14 9.241569
Rin27_15 in27_14 in27_15 9.241569
Rin27_16 in27_15 in27_16 9.241569
Rin27_17 in27_16 in27_17 9.241569
Rin27_18 in27_17 in27_18 9.241569
Rin27_19 in27_18 in27_19 9.241569
Rin27_20 in27_19 in27_20 9.241569
Rin27_21 in27_20 in27_21 9.241569
Rin27_22 in27_21 in27_22 9.241569
Rin27_23 in27_22 in27_23 9.241569
Rin27_24 in27_23 in27_24 9.241569
Rin27_25 in27_24 in27_25 9.241569
Rin27_26 in27_25 in27_26 9.241569
Rin27_27 in27_26 in27_27 9.241569
Rin27_28 in27_27 in27_28 9.241569
Rin27_29 in27 in27_29 9.241569
Rin27_30 in27_29 in27_30 9.241569
Rin27_31 in27_30 in27_31 9.241569
Rin27_32 in27_31 in27_32 9.241569
Rin27_33 in27_32 in27_33 9.241569
Rin27_34 in27_33 in27_34 9.241569
Rin27_35 in27_34 in27_35 9.241569
Rin27_36 in27_35 in27_36 9.241569
Rin27_37 in27_36 in27_37 9.241569
Rin27_38 in27_37 in27_38 9.241569
Rin27_39 in27_38 in27_39 9.241569
Rin27_40 in27_39 in27_40 9.241569
Rin27_41 in27_40 in27_41 9.241569
Rin27_42 in27_41 in27_42 9.241569
Rin27_43 in27_42 in27_43 9.241569
Rin27_44 in27_43 in27_44 9.241569
Rin27_45 in27_44 in27_45 9.241569
Rin27_46 in27_45 in27_46 9.241569
Rin27_47 in27_46 in27_47 9.241569
Rin27_48 in27_47 in27_48 9.241569
Rin27_49 in27_48 in27_49 9.241569
Rin27_50 in27_49 in27_50 9.241569
Rin27_51 in27_50 in27_51 9.241569
Rin27_52 in27_51 in27_52 9.241569
Rin27_53 in27_52 in27_53 9.241569
Rin27_54 in27_53 in27_54 9.241569
Rin27_55 in27_54 in27_55 9.241569
Rin27_56 in27_55 in27_56 9.241569
Rin27_57 in27 in27_57 9.241569
Rin27_58 in27_57 in27_58 9.241569
Rin27_59 in27_58 in27_59 9.241569
Rin27_60 in27_59 in27_60 9.241569
Rin27_61 in27_60 in27_61 9.241569
Rin27_62 in27_61 in27_62 9.241569
Rin27_63 in27_62 in27_63 9.241569
Rin27_64 in27_63 in27_64 9.241569
Rin27_65 in27_64 in27_65 9.241569
Rin27_66 in27_65 in27_66 9.241569
Rin27_67 in27_66 in27_67 9.241569
Rin27_68 in27_67 in27_68 9.241569
Rin27_69 in27_68 in27_69 9.241569
Rin27_70 in27_69 in27_70 9.241569
Rin27_71 in27_70 in27_71 9.241569
Rin27_72 in27_71 in27_72 9.241569
Rin27_73 in27_72 in27_73 9.241569
Rin27_74 in27_73 in27_74 9.241569
Rin27_75 in27_74 in27_75 9.241569
Rin27_76 in27_75 in27_76 9.241569
Rin27_77 in27_76 in27_77 9.241569
Rin27_78 in27_77 in27_78 9.241569
Rin27_79 in27_78 in27_79 9.241569
Rin27_80 in27_79 in27_80 9.241569
Rin27_81 in27_80 in27_81 9.241569
Rin27_82 in27_81 in27_82 9.241569
Rin27_83 in27_82 in27_83 9.241569
Rin27_84 in27_83 in27_84 9.241569
Rin28_1 in28 in28_1 9.241569
Rin28_2 in28_1 in28_2 9.241569
Rin28_3 in28_2 in28_3 9.241569
Rin28_4 in28_3 in28_4 9.241569
Rin28_5 in28_4 in28_5 9.241569
Rin28_6 in28_5 in28_6 9.241569
Rin28_7 in28_6 in28_7 9.241569
Rin28_8 in28_7 in28_8 9.241569
Rin28_9 in28_8 in28_9 9.241569
Rin28_10 in28_9 in28_10 9.241569
Rin28_11 in28_10 in28_11 9.241569
Rin28_12 in28_11 in28_12 9.241569
Rin28_13 in28_12 in28_13 9.241569
Rin28_14 in28_13 in28_14 9.241569
Rin28_15 in28_14 in28_15 9.241569
Rin28_16 in28_15 in28_16 9.241569
Rin28_17 in28_16 in28_17 9.241569
Rin28_18 in28_17 in28_18 9.241569
Rin28_19 in28_18 in28_19 9.241569
Rin28_20 in28_19 in28_20 9.241569
Rin28_21 in28_20 in28_21 9.241569
Rin28_22 in28_21 in28_22 9.241569
Rin28_23 in28_22 in28_23 9.241569
Rin28_24 in28_23 in28_24 9.241569
Rin28_25 in28_24 in28_25 9.241569
Rin28_26 in28_25 in28_26 9.241569
Rin28_27 in28_26 in28_27 9.241569
Rin28_28 in28_27 in28_28 9.241569
Rin28_29 in28 in28_29 9.241569
Rin28_30 in28_29 in28_30 9.241569
Rin28_31 in28_30 in28_31 9.241569
Rin28_32 in28_31 in28_32 9.241569
Rin28_33 in28_32 in28_33 9.241569
Rin28_34 in28_33 in28_34 9.241569
Rin28_35 in28_34 in28_35 9.241569
Rin28_36 in28_35 in28_36 9.241569
Rin28_37 in28_36 in28_37 9.241569
Rin28_38 in28_37 in28_38 9.241569
Rin28_39 in28_38 in28_39 9.241569
Rin28_40 in28_39 in28_40 9.241569
Rin28_41 in28_40 in28_41 9.241569
Rin28_42 in28_41 in28_42 9.241569
Rin28_43 in28_42 in28_43 9.241569
Rin28_44 in28_43 in28_44 9.241569
Rin28_45 in28_44 in28_45 9.241569
Rin28_46 in28_45 in28_46 9.241569
Rin28_47 in28_46 in28_47 9.241569
Rin28_48 in28_47 in28_48 9.241569
Rin28_49 in28_48 in28_49 9.241569
Rin28_50 in28_49 in28_50 9.241569
Rin28_51 in28_50 in28_51 9.241569
Rin28_52 in28_51 in28_52 9.241569
Rin28_53 in28_52 in28_53 9.241569
Rin28_54 in28_53 in28_54 9.241569
Rin28_55 in28_54 in28_55 9.241569
Rin28_56 in28_55 in28_56 9.241569
Rin28_57 in28 in28_57 9.241569
Rin28_58 in28_57 in28_58 9.241569
Rin28_59 in28_58 in28_59 9.241569
Rin28_60 in28_59 in28_60 9.241569
Rin28_61 in28_60 in28_61 9.241569
Rin28_62 in28_61 in28_62 9.241569
Rin28_63 in28_62 in28_63 9.241569
Rin28_64 in28_63 in28_64 9.241569
Rin28_65 in28_64 in28_65 9.241569
Rin28_66 in28_65 in28_66 9.241569
Rin28_67 in28_66 in28_67 9.241569
Rin28_68 in28_67 in28_68 9.241569
Rin28_69 in28_68 in28_69 9.241569
Rin28_70 in28_69 in28_70 9.241569
Rin28_71 in28_70 in28_71 9.241569
Rin28_72 in28_71 in28_72 9.241569
Rin28_73 in28_72 in28_73 9.241569
Rin28_74 in28_73 in28_74 9.241569
Rin28_75 in28_74 in28_75 9.241569
Rin28_76 in28_75 in28_76 9.241569
Rin28_77 in28_76 in28_77 9.241569
Rin28_78 in28_77 in28_78 9.241569
Rin28_79 in28_78 in28_79 9.241569
Rin28_80 in28_79 in28_80 9.241569
Rin28_81 in28_80 in28_81 9.241569
Rin28_82 in28_81 in28_82 9.241569
Rin28_83 in28_82 in28_83 9.241569
Rin28_84 in28_83 in28_84 9.241569
Rin29_1 in29 in29_1 9.241569
Rin29_2 in29_1 in29_2 9.241569
Rin29_3 in29_2 in29_3 9.241569
Rin29_4 in29_3 in29_4 9.241569
Rin29_5 in29_4 in29_5 9.241569
Rin29_6 in29_5 in29_6 9.241569
Rin29_7 in29_6 in29_7 9.241569
Rin29_8 in29_7 in29_8 9.241569
Rin29_9 in29_8 in29_9 9.241569
Rin29_10 in29_9 in29_10 9.241569
Rin29_11 in29_10 in29_11 9.241569
Rin29_12 in29_11 in29_12 9.241569
Rin29_13 in29_12 in29_13 9.241569
Rin29_14 in29_13 in29_14 9.241569
Rin29_15 in29_14 in29_15 9.241569
Rin29_16 in29_15 in29_16 9.241569
Rin29_17 in29_16 in29_17 9.241569
Rin29_18 in29_17 in29_18 9.241569
Rin29_19 in29_18 in29_19 9.241569
Rin29_20 in29_19 in29_20 9.241569
Rin29_21 in29_20 in29_21 9.241569
Rin29_22 in29_21 in29_22 9.241569
Rin29_23 in29_22 in29_23 9.241569
Rin29_24 in29_23 in29_24 9.241569
Rin29_25 in29_24 in29_25 9.241569
Rin29_26 in29_25 in29_26 9.241569
Rin29_27 in29_26 in29_27 9.241569
Rin29_28 in29_27 in29_28 9.241569
Rin29_29 in29 in29_29 9.241569
Rin29_30 in29_29 in29_30 9.241569
Rin29_31 in29_30 in29_31 9.241569
Rin29_32 in29_31 in29_32 9.241569
Rin29_33 in29_32 in29_33 9.241569
Rin29_34 in29_33 in29_34 9.241569
Rin29_35 in29_34 in29_35 9.241569
Rin29_36 in29_35 in29_36 9.241569
Rin29_37 in29_36 in29_37 9.241569
Rin29_38 in29_37 in29_38 9.241569
Rin29_39 in29_38 in29_39 9.241569
Rin29_40 in29_39 in29_40 9.241569
Rin29_41 in29_40 in29_41 9.241569
Rin29_42 in29_41 in29_42 9.241569
Rin29_43 in29_42 in29_43 9.241569
Rin29_44 in29_43 in29_44 9.241569
Rin29_45 in29_44 in29_45 9.241569
Rin29_46 in29_45 in29_46 9.241569
Rin29_47 in29_46 in29_47 9.241569
Rin29_48 in29_47 in29_48 9.241569
Rin29_49 in29_48 in29_49 9.241569
Rin29_50 in29_49 in29_50 9.241569
Rin29_51 in29_50 in29_51 9.241569
Rin29_52 in29_51 in29_52 9.241569
Rin29_53 in29_52 in29_53 9.241569
Rin29_54 in29_53 in29_54 9.241569
Rin29_55 in29_54 in29_55 9.241569
Rin29_56 in29_55 in29_56 9.241569
Rin29_57 in29 in29_57 9.241569
Rin29_58 in29_57 in29_58 9.241569
Rin29_59 in29_58 in29_59 9.241569
Rin29_60 in29_59 in29_60 9.241569
Rin29_61 in29_60 in29_61 9.241569
Rin29_62 in29_61 in29_62 9.241569
Rin29_63 in29_62 in29_63 9.241569
Rin29_64 in29_63 in29_64 9.241569
Rin29_65 in29_64 in29_65 9.241569
Rin29_66 in29_65 in29_66 9.241569
Rin29_67 in29_66 in29_67 9.241569
Rin29_68 in29_67 in29_68 9.241569
Rin29_69 in29_68 in29_69 9.241569
Rin29_70 in29_69 in29_70 9.241569
Rin29_71 in29_70 in29_71 9.241569
Rin29_72 in29_71 in29_72 9.241569
Rin29_73 in29_72 in29_73 9.241569
Rin29_74 in29_73 in29_74 9.241569
Rin29_75 in29_74 in29_75 9.241569
Rin29_76 in29_75 in29_76 9.241569
Rin29_77 in29_76 in29_77 9.241569
Rin29_78 in29_77 in29_78 9.241569
Rin29_79 in29_78 in29_79 9.241569
Rin29_80 in29_79 in29_80 9.241569
Rin29_81 in29_80 in29_81 9.241569
Rin29_82 in29_81 in29_82 9.241569
Rin29_83 in29_82 in29_83 9.241569
Rin29_84 in29_83 in29_84 9.241569
Rin30_1 in30 in30_1 9.241569
Rin30_2 in30_1 in30_2 9.241569
Rin30_3 in30_2 in30_3 9.241569
Rin30_4 in30_3 in30_4 9.241569
Rin30_5 in30_4 in30_5 9.241569
Rin30_6 in30_5 in30_6 9.241569
Rin30_7 in30_6 in30_7 9.241569
Rin30_8 in30_7 in30_8 9.241569
Rin30_9 in30_8 in30_9 9.241569
Rin30_10 in30_9 in30_10 9.241569
Rin30_11 in30_10 in30_11 9.241569
Rin30_12 in30_11 in30_12 9.241569
Rin30_13 in30_12 in30_13 9.241569
Rin30_14 in30_13 in30_14 9.241569
Rin30_15 in30_14 in30_15 9.241569
Rin30_16 in30_15 in30_16 9.241569
Rin30_17 in30_16 in30_17 9.241569
Rin30_18 in30_17 in30_18 9.241569
Rin30_19 in30_18 in30_19 9.241569
Rin30_20 in30_19 in30_20 9.241569
Rin30_21 in30_20 in30_21 9.241569
Rin30_22 in30_21 in30_22 9.241569
Rin30_23 in30_22 in30_23 9.241569
Rin30_24 in30_23 in30_24 9.241569
Rin30_25 in30_24 in30_25 9.241569
Rin30_26 in30_25 in30_26 9.241569
Rin30_27 in30_26 in30_27 9.241569
Rin30_28 in30_27 in30_28 9.241569
Rin30_29 in30 in30_29 9.241569
Rin30_30 in30_29 in30_30 9.241569
Rin30_31 in30_30 in30_31 9.241569
Rin30_32 in30_31 in30_32 9.241569
Rin30_33 in30_32 in30_33 9.241569
Rin30_34 in30_33 in30_34 9.241569
Rin30_35 in30_34 in30_35 9.241569
Rin30_36 in30_35 in30_36 9.241569
Rin30_37 in30_36 in30_37 9.241569
Rin30_38 in30_37 in30_38 9.241569
Rin30_39 in30_38 in30_39 9.241569
Rin30_40 in30_39 in30_40 9.241569
Rin30_41 in30_40 in30_41 9.241569
Rin30_42 in30_41 in30_42 9.241569
Rin30_43 in30_42 in30_43 9.241569
Rin30_44 in30_43 in30_44 9.241569
Rin30_45 in30_44 in30_45 9.241569
Rin30_46 in30_45 in30_46 9.241569
Rin30_47 in30_46 in30_47 9.241569
Rin30_48 in30_47 in30_48 9.241569
Rin30_49 in30_48 in30_49 9.241569
Rin30_50 in30_49 in30_50 9.241569
Rin30_51 in30_50 in30_51 9.241569
Rin30_52 in30_51 in30_52 9.241569
Rin30_53 in30_52 in30_53 9.241569
Rin30_54 in30_53 in30_54 9.241569
Rin30_55 in30_54 in30_55 9.241569
Rin30_56 in30_55 in30_56 9.241569
Rin30_57 in30 in30_57 9.241569
Rin30_58 in30_57 in30_58 9.241569
Rin30_59 in30_58 in30_59 9.241569
Rin30_60 in30_59 in30_60 9.241569
Rin30_61 in30_60 in30_61 9.241569
Rin30_62 in30_61 in30_62 9.241569
Rin30_63 in30_62 in30_63 9.241569
Rin30_64 in30_63 in30_64 9.241569
Rin30_65 in30_64 in30_65 9.241569
Rin30_66 in30_65 in30_66 9.241569
Rin30_67 in30_66 in30_67 9.241569
Rin30_68 in30_67 in30_68 9.241569
Rin30_69 in30_68 in30_69 9.241569
Rin30_70 in30_69 in30_70 9.241569
Rin30_71 in30_70 in30_71 9.241569
Rin30_72 in30_71 in30_72 9.241569
Rin30_73 in30_72 in30_73 9.241569
Rin30_74 in30_73 in30_74 9.241569
Rin30_75 in30_74 in30_75 9.241569
Rin30_76 in30_75 in30_76 9.241569
Rin30_77 in30_76 in30_77 9.241569
Rin30_78 in30_77 in30_78 9.241569
Rin30_79 in30_78 in30_79 9.241569
Rin30_80 in30_79 in30_80 9.241569
Rin30_81 in30_80 in30_81 9.241569
Rin30_82 in30_81 in30_82 9.241569
Rin30_83 in30_82 in30_83 9.241569
Rin30_84 in30_83 in30_84 9.241569
Rin31_1 in31 in31_1 9.241569
Rin31_2 in31_1 in31_2 9.241569
Rin31_3 in31_2 in31_3 9.241569
Rin31_4 in31_3 in31_4 9.241569
Rin31_5 in31_4 in31_5 9.241569
Rin31_6 in31_5 in31_6 9.241569
Rin31_7 in31_6 in31_7 9.241569
Rin31_8 in31_7 in31_8 9.241569
Rin31_9 in31_8 in31_9 9.241569
Rin31_10 in31_9 in31_10 9.241569
Rin31_11 in31_10 in31_11 9.241569
Rin31_12 in31_11 in31_12 9.241569
Rin31_13 in31_12 in31_13 9.241569
Rin31_14 in31_13 in31_14 9.241569
Rin31_15 in31_14 in31_15 9.241569
Rin31_16 in31_15 in31_16 9.241569
Rin31_17 in31_16 in31_17 9.241569
Rin31_18 in31_17 in31_18 9.241569
Rin31_19 in31_18 in31_19 9.241569
Rin31_20 in31_19 in31_20 9.241569
Rin31_21 in31_20 in31_21 9.241569
Rin31_22 in31_21 in31_22 9.241569
Rin31_23 in31_22 in31_23 9.241569
Rin31_24 in31_23 in31_24 9.241569
Rin31_25 in31_24 in31_25 9.241569
Rin31_26 in31_25 in31_26 9.241569
Rin31_27 in31_26 in31_27 9.241569
Rin31_28 in31_27 in31_28 9.241569
Rin31_29 in31 in31_29 9.241569
Rin31_30 in31_29 in31_30 9.241569
Rin31_31 in31_30 in31_31 9.241569
Rin31_32 in31_31 in31_32 9.241569
Rin31_33 in31_32 in31_33 9.241569
Rin31_34 in31_33 in31_34 9.241569
Rin31_35 in31_34 in31_35 9.241569
Rin31_36 in31_35 in31_36 9.241569
Rin31_37 in31_36 in31_37 9.241569
Rin31_38 in31_37 in31_38 9.241569
Rin31_39 in31_38 in31_39 9.241569
Rin31_40 in31_39 in31_40 9.241569
Rin31_41 in31_40 in31_41 9.241569
Rin31_42 in31_41 in31_42 9.241569
Rin31_43 in31_42 in31_43 9.241569
Rin31_44 in31_43 in31_44 9.241569
Rin31_45 in31_44 in31_45 9.241569
Rin31_46 in31_45 in31_46 9.241569
Rin31_47 in31_46 in31_47 9.241569
Rin31_48 in31_47 in31_48 9.241569
Rin31_49 in31_48 in31_49 9.241569
Rin31_50 in31_49 in31_50 9.241569
Rin31_51 in31_50 in31_51 9.241569
Rin31_52 in31_51 in31_52 9.241569
Rin31_53 in31_52 in31_53 9.241569
Rin31_54 in31_53 in31_54 9.241569
Rin31_55 in31_54 in31_55 9.241569
Rin31_56 in31_55 in31_56 9.241569
Rin31_57 in31 in31_57 9.241569
Rin31_58 in31_57 in31_58 9.241569
Rin31_59 in31_58 in31_59 9.241569
Rin31_60 in31_59 in31_60 9.241569
Rin31_61 in31_60 in31_61 9.241569
Rin31_62 in31_61 in31_62 9.241569
Rin31_63 in31_62 in31_63 9.241569
Rin31_64 in31_63 in31_64 9.241569
Rin31_65 in31_64 in31_65 9.241569
Rin31_66 in31_65 in31_66 9.241569
Rin31_67 in31_66 in31_67 9.241569
Rin31_68 in31_67 in31_68 9.241569
Rin31_69 in31_68 in31_69 9.241569
Rin31_70 in31_69 in31_70 9.241569
Rin31_71 in31_70 in31_71 9.241569
Rin31_72 in31_71 in31_72 9.241569
Rin31_73 in31_72 in31_73 9.241569
Rin31_74 in31_73 in31_74 9.241569
Rin31_75 in31_74 in31_75 9.241569
Rin31_76 in31_75 in31_76 9.241569
Rin31_77 in31_76 in31_77 9.241569
Rin31_78 in31_77 in31_78 9.241569
Rin31_79 in31_78 in31_79 9.241569
Rin31_80 in31_79 in31_80 9.241569
Rin31_81 in31_80 in31_81 9.241569
Rin31_82 in31_81 in31_82 9.241569
Rin31_83 in31_82 in31_83 9.241569
Rin31_84 in31_83 in31_84 9.241569
Rin32_1 in32 in32_1 9.241569
Rin32_2 in32_1 in32_2 9.241569
Rin32_3 in32_2 in32_3 9.241569
Rin32_4 in32_3 in32_4 9.241569
Rin32_5 in32_4 in32_5 9.241569
Rin32_6 in32_5 in32_6 9.241569
Rin32_7 in32_6 in32_7 9.241569
Rin32_8 in32_7 in32_8 9.241569
Rin32_9 in32_8 in32_9 9.241569
Rin32_10 in32_9 in32_10 9.241569
Rin32_11 in32_10 in32_11 9.241569
Rin32_12 in32_11 in32_12 9.241569
Rin32_13 in32_12 in32_13 9.241569
Rin32_14 in32_13 in32_14 9.241569
Rin32_15 in32_14 in32_15 9.241569
Rin32_16 in32_15 in32_16 9.241569
Rin32_17 in32_16 in32_17 9.241569
Rin32_18 in32_17 in32_18 9.241569
Rin32_19 in32_18 in32_19 9.241569
Rin32_20 in32_19 in32_20 9.241569
Rin32_21 in32_20 in32_21 9.241569
Rin32_22 in32_21 in32_22 9.241569
Rin32_23 in32_22 in32_23 9.241569
Rin32_24 in32_23 in32_24 9.241569
Rin32_25 in32_24 in32_25 9.241569
Rin32_26 in32_25 in32_26 9.241569
Rin32_27 in32_26 in32_27 9.241569
Rin32_28 in32_27 in32_28 9.241569
Rin32_29 in32 in32_29 9.241569
Rin32_30 in32_29 in32_30 9.241569
Rin32_31 in32_30 in32_31 9.241569
Rin32_32 in32_31 in32_32 9.241569
Rin32_33 in32_32 in32_33 9.241569
Rin32_34 in32_33 in32_34 9.241569
Rin32_35 in32_34 in32_35 9.241569
Rin32_36 in32_35 in32_36 9.241569
Rin32_37 in32_36 in32_37 9.241569
Rin32_38 in32_37 in32_38 9.241569
Rin32_39 in32_38 in32_39 9.241569
Rin32_40 in32_39 in32_40 9.241569
Rin32_41 in32_40 in32_41 9.241569
Rin32_42 in32_41 in32_42 9.241569
Rin32_43 in32_42 in32_43 9.241569
Rin32_44 in32_43 in32_44 9.241569
Rin32_45 in32_44 in32_45 9.241569
Rin32_46 in32_45 in32_46 9.241569
Rin32_47 in32_46 in32_47 9.241569
Rin32_48 in32_47 in32_48 9.241569
Rin32_49 in32_48 in32_49 9.241569
Rin32_50 in32_49 in32_50 9.241569
Rin32_51 in32_50 in32_51 9.241569
Rin32_52 in32_51 in32_52 9.241569
Rin32_53 in32_52 in32_53 9.241569
Rin32_54 in32_53 in32_54 9.241569
Rin32_55 in32_54 in32_55 9.241569
Rin32_56 in32_55 in32_56 9.241569
Rin32_57 in32 in32_57 9.241569
Rin32_58 in32_57 in32_58 9.241569
Rin32_59 in32_58 in32_59 9.241569
Rin32_60 in32_59 in32_60 9.241569
Rin32_61 in32_60 in32_61 9.241569
Rin32_62 in32_61 in32_62 9.241569
Rin32_63 in32_62 in32_63 9.241569
Rin32_64 in32_63 in32_64 9.241569
Rin32_65 in32_64 in32_65 9.241569
Rin32_66 in32_65 in32_66 9.241569
Rin32_67 in32_66 in32_67 9.241569
Rin32_68 in32_67 in32_68 9.241569
Rin32_69 in32_68 in32_69 9.241569
Rin32_70 in32_69 in32_70 9.241569
Rin32_71 in32_70 in32_71 9.241569
Rin32_72 in32_71 in32_72 9.241569
Rin32_73 in32_72 in32_73 9.241569
Rin32_74 in32_73 in32_74 9.241569
Rin32_75 in32_74 in32_75 9.241569
Rin32_76 in32_75 in32_76 9.241569
Rin32_77 in32_76 in32_77 9.241569
Rin32_78 in32_77 in32_78 9.241569
Rin32_79 in32_78 in32_79 9.241569
Rin32_80 in32_79 in32_80 9.241569
Rin32_81 in32_80 in32_81 9.241569
Rin32_82 in32_81 in32_82 9.241569
Rin32_83 in32_82 in32_83 9.241569
Rin32_84 in32_83 in32_84 9.241569
Rin33_1 in33 in33_1 9.241569
Rin33_2 in33_1 in33_2 9.241569
Rin33_3 in33_2 in33_3 9.241569
Rin33_4 in33_3 in33_4 9.241569
Rin33_5 in33_4 in33_5 9.241569
Rin33_6 in33_5 in33_6 9.241569
Rin33_7 in33_6 in33_7 9.241569
Rin33_8 in33_7 in33_8 9.241569
Rin33_9 in33_8 in33_9 9.241569
Rin33_10 in33_9 in33_10 9.241569
Rin33_11 in33_10 in33_11 9.241569
Rin33_12 in33_11 in33_12 9.241569
Rin33_13 in33_12 in33_13 9.241569
Rin33_14 in33_13 in33_14 9.241569
Rin33_15 in33_14 in33_15 9.241569
Rin33_16 in33_15 in33_16 9.241569
Rin33_17 in33_16 in33_17 9.241569
Rin33_18 in33_17 in33_18 9.241569
Rin33_19 in33_18 in33_19 9.241569
Rin33_20 in33_19 in33_20 9.241569
Rin33_21 in33_20 in33_21 9.241569
Rin33_22 in33_21 in33_22 9.241569
Rin33_23 in33_22 in33_23 9.241569
Rin33_24 in33_23 in33_24 9.241569
Rin33_25 in33_24 in33_25 9.241569
Rin33_26 in33_25 in33_26 9.241569
Rin33_27 in33_26 in33_27 9.241569
Rin33_28 in33_27 in33_28 9.241569
Rin33_29 in33 in33_29 9.241569
Rin33_30 in33_29 in33_30 9.241569
Rin33_31 in33_30 in33_31 9.241569
Rin33_32 in33_31 in33_32 9.241569
Rin33_33 in33_32 in33_33 9.241569
Rin33_34 in33_33 in33_34 9.241569
Rin33_35 in33_34 in33_35 9.241569
Rin33_36 in33_35 in33_36 9.241569
Rin33_37 in33_36 in33_37 9.241569
Rin33_38 in33_37 in33_38 9.241569
Rin33_39 in33_38 in33_39 9.241569
Rin33_40 in33_39 in33_40 9.241569
Rin33_41 in33_40 in33_41 9.241569
Rin33_42 in33_41 in33_42 9.241569
Rin33_43 in33_42 in33_43 9.241569
Rin33_44 in33_43 in33_44 9.241569
Rin33_45 in33_44 in33_45 9.241569
Rin33_46 in33_45 in33_46 9.241569
Rin33_47 in33_46 in33_47 9.241569
Rin33_48 in33_47 in33_48 9.241569
Rin33_49 in33_48 in33_49 9.241569
Rin33_50 in33_49 in33_50 9.241569
Rin33_51 in33_50 in33_51 9.241569
Rin33_52 in33_51 in33_52 9.241569
Rin33_53 in33_52 in33_53 9.241569
Rin33_54 in33_53 in33_54 9.241569
Rin33_55 in33_54 in33_55 9.241569
Rin33_56 in33_55 in33_56 9.241569
Rin33_57 in33 in33_57 9.241569
Rin33_58 in33_57 in33_58 9.241569
Rin33_59 in33_58 in33_59 9.241569
Rin33_60 in33_59 in33_60 9.241569
Rin33_61 in33_60 in33_61 9.241569
Rin33_62 in33_61 in33_62 9.241569
Rin33_63 in33_62 in33_63 9.241569
Rin33_64 in33_63 in33_64 9.241569
Rin33_65 in33_64 in33_65 9.241569
Rin33_66 in33_65 in33_66 9.241569
Rin33_67 in33_66 in33_67 9.241569
Rin33_68 in33_67 in33_68 9.241569
Rin33_69 in33_68 in33_69 9.241569
Rin33_70 in33_69 in33_70 9.241569
Rin33_71 in33_70 in33_71 9.241569
Rin33_72 in33_71 in33_72 9.241569
Rin33_73 in33_72 in33_73 9.241569
Rin33_74 in33_73 in33_74 9.241569
Rin33_75 in33_74 in33_75 9.241569
Rin33_76 in33_75 in33_76 9.241569
Rin33_77 in33_76 in33_77 9.241569
Rin33_78 in33_77 in33_78 9.241569
Rin33_79 in33_78 in33_79 9.241569
Rin33_80 in33_79 in33_80 9.241569
Rin33_81 in33_80 in33_81 9.241569
Rin33_82 in33_81 in33_82 9.241569
Rin33_83 in33_82 in33_83 9.241569
Rin33_84 in33_83 in33_84 9.241569
Rin34_1 in34 in34_1 9.241569
Rin34_2 in34_1 in34_2 9.241569
Rin34_3 in34_2 in34_3 9.241569
Rin34_4 in34_3 in34_4 9.241569
Rin34_5 in34_4 in34_5 9.241569
Rin34_6 in34_5 in34_6 9.241569
Rin34_7 in34_6 in34_7 9.241569
Rin34_8 in34_7 in34_8 9.241569
Rin34_9 in34_8 in34_9 9.241569
Rin34_10 in34_9 in34_10 9.241569
Rin34_11 in34_10 in34_11 9.241569
Rin34_12 in34_11 in34_12 9.241569
Rin34_13 in34_12 in34_13 9.241569
Rin34_14 in34_13 in34_14 9.241569
Rin34_15 in34_14 in34_15 9.241569
Rin34_16 in34_15 in34_16 9.241569
Rin34_17 in34_16 in34_17 9.241569
Rin34_18 in34_17 in34_18 9.241569
Rin34_19 in34_18 in34_19 9.241569
Rin34_20 in34_19 in34_20 9.241569
Rin34_21 in34_20 in34_21 9.241569
Rin34_22 in34_21 in34_22 9.241569
Rin34_23 in34_22 in34_23 9.241569
Rin34_24 in34_23 in34_24 9.241569
Rin34_25 in34_24 in34_25 9.241569
Rin34_26 in34_25 in34_26 9.241569
Rin34_27 in34_26 in34_27 9.241569
Rin34_28 in34_27 in34_28 9.241569
Rin34_29 in34 in34_29 9.241569
Rin34_30 in34_29 in34_30 9.241569
Rin34_31 in34_30 in34_31 9.241569
Rin34_32 in34_31 in34_32 9.241569
Rin34_33 in34_32 in34_33 9.241569
Rin34_34 in34_33 in34_34 9.241569
Rin34_35 in34_34 in34_35 9.241569
Rin34_36 in34_35 in34_36 9.241569
Rin34_37 in34_36 in34_37 9.241569
Rin34_38 in34_37 in34_38 9.241569
Rin34_39 in34_38 in34_39 9.241569
Rin34_40 in34_39 in34_40 9.241569
Rin34_41 in34_40 in34_41 9.241569
Rin34_42 in34_41 in34_42 9.241569
Rin34_43 in34_42 in34_43 9.241569
Rin34_44 in34_43 in34_44 9.241569
Rin34_45 in34_44 in34_45 9.241569
Rin34_46 in34_45 in34_46 9.241569
Rin34_47 in34_46 in34_47 9.241569
Rin34_48 in34_47 in34_48 9.241569
Rin34_49 in34_48 in34_49 9.241569
Rin34_50 in34_49 in34_50 9.241569
Rin34_51 in34_50 in34_51 9.241569
Rin34_52 in34_51 in34_52 9.241569
Rin34_53 in34_52 in34_53 9.241569
Rin34_54 in34_53 in34_54 9.241569
Rin34_55 in34_54 in34_55 9.241569
Rin34_56 in34_55 in34_56 9.241569
Rin34_57 in34 in34_57 9.241569
Rin34_58 in34_57 in34_58 9.241569
Rin34_59 in34_58 in34_59 9.241569
Rin34_60 in34_59 in34_60 9.241569
Rin34_61 in34_60 in34_61 9.241569
Rin34_62 in34_61 in34_62 9.241569
Rin34_63 in34_62 in34_63 9.241569
Rin34_64 in34_63 in34_64 9.241569
Rin34_65 in34_64 in34_65 9.241569
Rin34_66 in34_65 in34_66 9.241569
Rin34_67 in34_66 in34_67 9.241569
Rin34_68 in34_67 in34_68 9.241569
Rin34_69 in34_68 in34_69 9.241569
Rin34_70 in34_69 in34_70 9.241569
Rin34_71 in34_70 in34_71 9.241569
Rin34_72 in34_71 in34_72 9.241569
Rin34_73 in34_72 in34_73 9.241569
Rin34_74 in34_73 in34_74 9.241569
Rin34_75 in34_74 in34_75 9.241569
Rin34_76 in34_75 in34_76 9.241569
Rin34_77 in34_76 in34_77 9.241569
Rin34_78 in34_77 in34_78 9.241569
Rin34_79 in34_78 in34_79 9.241569
Rin34_80 in34_79 in34_80 9.241569
Rin34_81 in34_80 in34_81 9.241569
Rin34_82 in34_81 in34_82 9.241569
Rin34_83 in34_82 in34_83 9.241569
Rin34_84 in34_83 in34_84 9.241569
Rin35_1 in35 in35_1 9.241569
Rin35_2 in35_1 in35_2 9.241569
Rin35_3 in35_2 in35_3 9.241569
Rin35_4 in35_3 in35_4 9.241569
Rin35_5 in35_4 in35_5 9.241569
Rin35_6 in35_5 in35_6 9.241569
Rin35_7 in35_6 in35_7 9.241569
Rin35_8 in35_7 in35_8 9.241569
Rin35_9 in35_8 in35_9 9.241569
Rin35_10 in35_9 in35_10 9.241569
Rin35_11 in35_10 in35_11 9.241569
Rin35_12 in35_11 in35_12 9.241569
Rin35_13 in35_12 in35_13 9.241569
Rin35_14 in35_13 in35_14 9.241569
Rin35_15 in35_14 in35_15 9.241569
Rin35_16 in35_15 in35_16 9.241569
Rin35_17 in35_16 in35_17 9.241569
Rin35_18 in35_17 in35_18 9.241569
Rin35_19 in35_18 in35_19 9.241569
Rin35_20 in35_19 in35_20 9.241569
Rin35_21 in35_20 in35_21 9.241569
Rin35_22 in35_21 in35_22 9.241569
Rin35_23 in35_22 in35_23 9.241569
Rin35_24 in35_23 in35_24 9.241569
Rin35_25 in35_24 in35_25 9.241569
Rin35_26 in35_25 in35_26 9.241569
Rin35_27 in35_26 in35_27 9.241569
Rin35_28 in35_27 in35_28 9.241569
Rin35_29 in35 in35_29 9.241569
Rin35_30 in35_29 in35_30 9.241569
Rin35_31 in35_30 in35_31 9.241569
Rin35_32 in35_31 in35_32 9.241569
Rin35_33 in35_32 in35_33 9.241569
Rin35_34 in35_33 in35_34 9.241569
Rin35_35 in35_34 in35_35 9.241569
Rin35_36 in35_35 in35_36 9.241569
Rin35_37 in35_36 in35_37 9.241569
Rin35_38 in35_37 in35_38 9.241569
Rin35_39 in35_38 in35_39 9.241569
Rin35_40 in35_39 in35_40 9.241569
Rin35_41 in35_40 in35_41 9.241569
Rin35_42 in35_41 in35_42 9.241569
Rin35_43 in35_42 in35_43 9.241569
Rin35_44 in35_43 in35_44 9.241569
Rin35_45 in35_44 in35_45 9.241569
Rin35_46 in35_45 in35_46 9.241569
Rin35_47 in35_46 in35_47 9.241569
Rin35_48 in35_47 in35_48 9.241569
Rin35_49 in35_48 in35_49 9.241569
Rin35_50 in35_49 in35_50 9.241569
Rin35_51 in35_50 in35_51 9.241569
Rin35_52 in35_51 in35_52 9.241569
Rin35_53 in35_52 in35_53 9.241569
Rin35_54 in35_53 in35_54 9.241569
Rin35_55 in35_54 in35_55 9.241569
Rin35_56 in35_55 in35_56 9.241569
Rin35_57 in35 in35_57 9.241569
Rin35_58 in35_57 in35_58 9.241569
Rin35_59 in35_58 in35_59 9.241569
Rin35_60 in35_59 in35_60 9.241569
Rin35_61 in35_60 in35_61 9.241569
Rin35_62 in35_61 in35_62 9.241569
Rin35_63 in35_62 in35_63 9.241569
Rin35_64 in35_63 in35_64 9.241569
Rin35_65 in35_64 in35_65 9.241569
Rin35_66 in35_65 in35_66 9.241569
Rin35_67 in35_66 in35_67 9.241569
Rin35_68 in35_67 in35_68 9.241569
Rin35_69 in35_68 in35_69 9.241569
Rin35_70 in35_69 in35_70 9.241569
Rin35_71 in35_70 in35_71 9.241569
Rin35_72 in35_71 in35_72 9.241569
Rin35_73 in35_72 in35_73 9.241569
Rin35_74 in35_73 in35_74 9.241569
Rin35_75 in35_74 in35_75 9.241569
Rin35_76 in35_75 in35_76 9.241569
Rin35_77 in35_76 in35_77 9.241569
Rin35_78 in35_77 in35_78 9.241569
Rin35_79 in35_78 in35_79 9.241569
Rin35_80 in35_79 in35_80 9.241569
Rin35_81 in35_80 in35_81 9.241569
Rin35_82 in35_81 in35_82 9.241569
Rin35_83 in35_82 in35_83 9.241569
Rin35_84 in35_83 in35_84 9.241569
Rin36_1 in36 in36_1 9.241569
Rin36_2 in36_1 in36_2 9.241569
Rin36_3 in36_2 in36_3 9.241569
Rin36_4 in36_3 in36_4 9.241569
Rin36_5 in36_4 in36_5 9.241569
Rin36_6 in36_5 in36_6 9.241569
Rin36_7 in36_6 in36_7 9.241569
Rin36_8 in36_7 in36_8 9.241569
Rin36_9 in36_8 in36_9 9.241569
Rin36_10 in36_9 in36_10 9.241569
Rin36_11 in36_10 in36_11 9.241569
Rin36_12 in36_11 in36_12 9.241569
Rin36_13 in36_12 in36_13 9.241569
Rin36_14 in36_13 in36_14 9.241569
Rin36_15 in36_14 in36_15 9.241569
Rin36_16 in36_15 in36_16 9.241569
Rin36_17 in36_16 in36_17 9.241569
Rin36_18 in36_17 in36_18 9.241569
Rin36_19 in36_18 in36_19 9.241569
Rin36_20 in36_19 in36_20 9.241569
Rin36_21 in36_20 in36_21 9.241569
Rin36_22 in36_21 in36_22 9.241569
Rin36_23 in36_22 in36_23 9.241569
Rin36_24 in36_23 in36_24 9.241569
Rin36_25 in36_24 in36_25 9.241569
Rin36_26 in36_25 in36_26 9.241569
Rin36_27 in36_26 in36_27 9.241569
Rin36_28 in36_27 in36_28 9.241569
Rin36_29 in36 in36_29 9.241569
Rin36_30 in36_29 in36_30 9.241569
Rin36_31 in36_30 in36_31 9.241569
Rin36_32 in36_31 in36_32 9.241569
Rin36_33 in36_32 in36_33 9.241569
Rin36_34 in36_33 in36_34 9.241569
Rin36_35 in36_34 in36_35 9.241569
Rin36_36 in36_35 in36_36 9.241569
Rin36_37 in36_36 in36_37 9.241569
Rin36_38 in36_37 in36_38 9.241569
Rin36_39 in36_38 in36_39 9.241569
Rin36_40 in36_39 in36_40 9.241569
Rin36_41 in36_40 in36_41 9.241569
Rin36_42 in36_41 in36_42 9.241569
Rin36_43 in36_42 in36_43 9.241569
Rin36_44 in36_43 in36_44 9.241569
Rin36_45 in36_44 in36_45 9.241569
Rin36_46 in36_45 in36_46 9.241569
Rin36_47 in36_46 in36_47 9.241569
Rin36_48 in36_47 in36_48 9.241569
Rin36_49 in36_48 in36_49 9.241569
Rin36_50 in36_49 in36_50 9.241569
Rin36_51 in36_50 in36_51 9.241569
Rin36_52 in36_51 in36_52 9.241569
Rin36_53 in36_52 in36_53 9.241569
Rin36_54 in36_53 in36_54 9.241569
Rin36_55 in36_54 in36_55 9.241569
Rin36_56 in36_55 in36_56 9.241569
Rin36_57 in36 in36_57 9.241569
Rin36_58 in36_57 in36_58 9.241569
Rin36_59 in36_58 in36_59 9.241569
Rin36_60 in36_59 in36_60 9.241569
Rin36_61 in36_60 in36_61 9.241569
Rin36_62 in36_61 in36_62 9.241569
Rin36_63 in36_62 in36_63 9.241569
Rin36_64 in36_63 in36_64 9.241569
Rin36_65 in36_64 in36_65 9.241569
Rin36_66 in36_65 in36_66 9.241569
Rin36_67 in36_66 in36_67 9.241569
Rin36_68 in36_67 in36_68 9.241569
Rin36_69 in36_68 in36_69 9.241569
Rin36_70 in36_69 in36_70 9.241569
Rin36_71 in36_70 in36_71 9.241569
Rin36_72 in36_71 in36_72 9.241569
Rin36_73 in36_72 in36_73 9.241569
Rin36_74 in36_73 in36_74 9.241569
Rin36_75 in36_74 in36_75 9.241569
Rin36_76 in36_75 in36_76 9.241569
Rin36_77 in36_76 in36_77 9.241569
Rin36_78 in36_77 in36_78 9.241569
Rin36_79 in36_78 in36_79 9.241569
Rin36_80 in36_79 in36_80 9.241569
Rin36_81 in36_80 in36_81 9.241569
Rin36_82 in36_81 in36_82 9.241569
Rin36_83 in36_82 in36_83 9.241569
Rin36_84 in36_83 in36_84 9.241569
Rin37_1 in37 in37_1 9.241569
Rin37_2 in37_1 in37_2 9.241569
Rin37_3 in37_2 in37_3 9.241569
Rin37_4 in37_3 in37_4 9.241569
Rin37_5 in37_4 in37_5 9.241569
Rin37_6 in37_5 in37_6 9.241569
Rin37_7 in37_6 in37_7 9.241569
Rin37_8 in37_7 in37_8 9.241569
Rin37_9 in37_8 in37_9 9.241569
Rin37_10 in37_9 in37_10 9.241569
Rin37_11 in37_10 in37_11 9.241569
Rin37_12 in37_11 in37_12 9.241569
Rin37_13 in37_12 in37_13 9.241569
Rin37_14 in37_13 in37_14 9.241569
Rin37_15 in37_14 in37_15 9.241569
Rin37_16 in37_15 in37_16 9.241569
Rin37_17 in37_16 in37_17 9.241569
Rin37_18 in37_17 in37_18 9.241569
Rin37_19 in37_18 in37_19 9.241569
Rin37_20 in37_19 in37_20 9.241569
Rin37_21 in37_20 in37_21 9.241569
Rin37_22 in37_21 in37_22 9.241569
Rin37_23 in37_22 in37_23 9.241569
Rin37_24 in37_23 in37_24 9.241569
Rin37_25 in37_24 in37_25 9.241569
Rin37_26 in37_25 in37_26 9.241569
Rin37_27 in37_26 in37_27 9.241569
Rin37_28 in37_27 in37_28 9.241569
Rin37_29 in37 in37_29 9.241569
Rin37_30 in37_29 in37_30 9.241569
Rin37_31 in37_30 in37_31 9.241569
Rin37_32 in37_31 in37_32 9.241569
Rin37_33 in37_32 in37_33 9.241569
Rin37_34 in37_33 in37_34 9.241569
Rin37_35 in37_34 in37_35 9.241569
Rin37_36 in37_35 in37_36 9.241569
Rin37_37 in37_36 in37_37 9.241569
Rin37_38 in37_37 in37_38 9.241569
Rin37_39 in37_38 in37_39 9.241569
Rin37_40 in37_39 in37_40 9.241569
Rin37_41 in37_40 in37_41 9.241569
Rin37_42 in37_41 in37_42 9.241569
Rin37_43 in37_42 in37_43 9.241569
Rin37_44 in37_43 in37_44 9.241569
Rin37_45 in37_44 in37_45 9.241569
Rin37_46 in37_45 in37_46 9.241569
Rin37_47 in37_46 in37_47 9.241569
Rin37_48 in37_47 in37_48 9.241569
Rin37_49 in37_48 in37_49 9.241569
Rin37_50 in37_49 in37_50 9.241569
Rin37_51 in37_50 in37_51 9.241569
Rin37_52 in37_51 in37_52 9.241569
Rin37_53 in37_52 in37_53 9.241569
Rin37_54 in37_53 in37_54 9.241569
Rin37_55 in37_54 in37_55 9.241569
Rin37_56 in37_55 in37_56 9.241569
Rin37_57 in37 in37_57 9.241569
Rin37_58 in37_57 in37_58 9.241569
Rin37_59 in37_58 in37_59 9.241569
Rin37_60 in37_59 in37_60 9.241569
Rin37_61 in37_60 in37_61 9.241569
Rin37_62 in37_61 in37_62 9.241569
Rin37_63 in37_62 in37_63 9.241569
Rin37_64 in37_63 in37_64 9.241569
Rin37_65 in37_64 in37_65 9.241569
Rin37_66 in37_65 in37_66 9.241569
Rin37_67 in37_66 in37_67 9.241569
Rin37_68 in37_67 in37_68 9.241569
Rin37_69 in37_68 in37_69 9.241569
Rin37_70 in37_69 in37_70 9.241569
Rin37_71 in37_70 in37_71 9.241569
Rin37_72 in37_71 in37_72 9.241569
Rin37_73 in37_72 in37_73 9.241569
Rin37_74 in37_73 in37_74 9.241569
Rin37_75 in37_74 in37_75 9.241569
Rin37_76 in37_75 in37_76 9.241569
Rin37_77 in37_76 in37_77 9.241569
Rin37_78 in37_77 in37_78 9.241569
Rin37_79 in37_78 in37_79 9.241569
Rin37_80 in37_79 in37_80 9.241569
Rin37_81 in37_80 in37_81 9.241569
Rin37_82 in37_81 in37_82 9.241569
Rin37_83 in37_82 in37_83 9.241569
Rin37_84 in37_83 in37_84 9.241569
Rin38_1 in38 in38_1 9.241569
Rin38_2 in38_1 in38_2 9.241569
Rin38_3 in38_2 in38_3 9.241569
Rin38_4 in38_3 in38_4 9.241569
Rin38_5 in38_4 in38_5 9.241569
Rin38_6 in38_5 in38_6 9.241569
Rin38_7 in38_6 in38_7 9.241569
Rin38_8 in38_7 in38_8 9.241569
Rin38_9 in38_8 in38_9 9.241569
Rin38_10 in38_9 in38_10 9.241569
Rin38_11 in38_10 in38_11 9.241569
Rin38_12 in38_11 in38_12 9.241569
Rin38_13 in38_12 in38_13 9.241569
Rin38_14 in38_13 in38_14 9.241569
Rin38_15 in38_14 in38_15 9.241569
Rin38_16 in38_15 in38_16 9.241569
Rin38_17 in38_16 in38_17 9.241569
Rin38_18 in38_17 in38_18 9.241569
Rin38_19 in38_18 in38_19 9.241569
Rin38_20 in38_19 in38_20 9.241569
Rin38_21 in38_20 in38_21 9.241569
Rin38_22 in38_21 in38_22 9.241569
Rin38_23 in38_22 in38_23 9.241569
Rin38_24 in38_23 in38_24 9.241569
Rin38_25 in38_24 in38_25 9.241569
Rin38_26 in38_25 in38_26 9.241569
Rin38_27 in38_26 in38_27 9.241569
Rin38_28 in38_27 in38_28 9.241569
Rin38_29 in38 in38_29 9.241569
Rin38_30 in38_29 in38_30 9.241569
Rin38_31 in38_30 in38_31 9.241569
Rin38_32 in38_31 in38_32 9.241569
Rin38_33 in38_32 in38_33 9.241569
Rin38_34 in38_33 in38_34 9.241569
Rin38_35 in38_34 in38_35 9.241569
Rin38_36 in38_35 in38_36 9.241569
Rin38_37 in38_36 in38_37 9.241569
Rin38_38 in38_37 in38_38 9.241569
Rin38_39 in38_38 in38_39 9.241569
Rin38_40 in38_39 in38_40 9.241569
Rin38_41 in38_40 in38_41 9.241569
Rin38_42 in38_41 in38_42 9.241569
Rin38_43 in38_42 in38_43 9.241569
Rin38_44 in38_43 in38_44 9.241569
Rin38_45 in38_44 in38_45 9.241569
Rin38_46 in38_45 in38_46 9.241569
Rin38_47 in38_46 in38_47 9.241569
Rin38_48 in38_47 in38_48 9.241569
Rin38_49 in38_48 in38_49 9.241569
Rin38_50 in38_49 in38_50 9.241569
Rin38_51 in38_50 in38_51 9.241569
Rin38_52 in38_51 in38_52 9.241569
Rin38_53 in38_52 in38_53 9.241569
Rin38_54 in38_53 in38_54 9.241569
Rin38_55 in38_54 in38_55 9.241569
Rin38_56 in38_55 in38_56 9.241569
Rin38_57 in38 in38_57 9.241569
Rin38_58 in38_57 in38_58 9.241569
Rin38_59 in38_58 in38_59 9.241569
Rin38_60 in38_59 in38_60 9.241569
Rin38_61 in38_60 in38_61 9.241569
Rin38_62 in38_61 in38_62 9.241569
Rin38_63 in38_62 in38_63 9.241569
Rin38_64 in38_63 in38_64 9.241569
Rin38_65 in38_64 in38_65 9.241569
Rin38_66 in38_65 in38_66 9.241569
Rin38_67 in38_66 in38_67 9.241569
Rin38_68 in38_67 in38_68 9.241569
Rin38_69 in38_68 in38_69 9.241569
Rin38_70 in38_69 in38_70 9.241569
Rin38_71 in38_70 in38_71 9.241569
Rin38_72 in38_71 in38_72 9.241569
Rin38_73 in38_72 in38_73 9.241569
Rin38_74 in38_73 in38_74 9.241569
Rin38_75 in38_74 in38_75 9.241569
Rin38_76 in38_75 in38_76 9.241569
Rin38_77 in38_76 in38_77 9.241569
Rin38_78 in38_77 in38_78 9.241569
Rin38_79 in38_78 in38_79 9.241569
Rin38_80 in38_79 in38_80 9.241569
Rin38_81 in38_80 in38_81 9.241569
Rin38_82 in38_81 in38_82 9.241569
Rin38_83 in38_82 in38_83 9.241569
Rin38_84 in38_83 in38_84 9.241569
Rin39_1 in39 in39_1 9.241569
Rin39_2 in39_1 in39_2 9.241569
Rin39_3 in39_2 in39_3 9.241569
Rin39_4 in39_3 in39_4 9.241569
Rin39_5 in39_4 in39_5 9.241569
Rin39_6 in39_5 in39_6 9.241569
Rin39_7 in39_6 in39_7 9.241569
Rin39_8 in39_7 in39_8 9.241569
Rin39_9 in39_8 in39_9 9.241569
Rin39_10 in39_9 in39_10 9.241569
Rin39_11 in39_10 in39_11 9.241569
Rin39_12 in39_11 in39_12 9.241569
Rin39_13 in39_12 in39_13 9.241569
Rin39_14 in39_13 in39_14 9.241569
Rin39_15 in39_14 in39_15 9.241569
Rin39_16 in39_15 in39_16 9.241569
Rin39_17 in39_16 in39_17 9.241569
Rin39_18 in39_17 in39_18 9.241569
Rin39_19 in39_18 in39_19 9.241569
Rin39_20 in39_19 in39_20 9.241569
Rin39_21 in39_20 in39_21 9.241569
Rin39_22 in39_21 in39_22 9.241569
Rin39_23 in39_22 in39_23 9.241569
Rin39_24 in39_23 in39_24 9.241569
Rin39_25 in39_24 in39_25 9.241569
Rin39_26 in39_25 in39_26 9.241569
Rin39_27 in39_26 in39_27 9.241569
Rin39_28 in39_27 in39_28 9.241569
Rin39_29 in39 in39_29 9.241569
Rin39_30 in39_29 in39_30 9.241569
Rin39_31 in39_30 in39_31 9.241569
Rin39_32 in39_31 in39_32 9.241569
Rin39_33 in39_32 in39_33 9.241569
Rin39_34 in39_33 in39_34 9.241569
Rin39_35 in39_34 in39_35 9.241569
Rin39_36 in39_35 in39_36 9.241569
Rin39_37 in39_36 in39_37 9.241569
Rin39_38 in39_37 in39_38 9.241569
Rin39_39 in39_38 in39_39 9.241569
Rin39_40 in39_39 in39_40 9.241569
Rin39_41 in39_40 in39_41 9.241569
Rin39_42 in39_41 in39_42 9.241569
Rin39_43 in39_42 in39_43 9.241569
Rin39_44 in39_43 in39_44 9.241569
Rin39_45 in39_44 in39_45 9.241569
Rin39_46 in39_45 in39_46 9.241569
Rin39_47 in39_46 in39_47 9.241569
Rin39_48 in39_47 in39_48 9.241569
Rin39_49 in39_48 in39_49 9.241569
Rin39_50 in39_49 in39_50 9.241569
Rin39_51 in39_50 in39_51 9.241569
Rin39_52 in39_51 in39_52 9.241569
Rin39_53 in39_52 in39_53 9.241569
Rin39_54 in39_53 in39_54 9.241569
Rin39_55 in39_54 in39_55 9.241569
Rin39_56 in39_55 in39_56 9.241569
Rin39_57 in39 in39_57 9.241569
Rin39_58 in39_57 in39_58 9.241569
Rin39_59 in39_58 in39_59 9.241569
Rin39_60 in39_59 in39_60 9.241569
Rin39_61 in39_60 in39_61 9.241569
Rin39_62 in39_61 in39_62 9.241569
Rin39_63 in39_62 in39_63 9.241569
Rin39_64 in39_63 in39_64 9.241569
Rin39_65 in39_64 in39_65 9.241569
Rin39_66 in39_65 in39_66 9.241569
Rin39_67 in39_66 in39_67 9.241569
Rin39_68 in39_67 in39_68 9.241569
Rin39_69 in39_68 in39_69 9.241569
Rin39_70 in39_69 in39_70 9.241569
Rin39_71 in39_70 in39_71 9.241569
Rin39_72 in39_71 in39_72 9.241569
Rin39_73 in39_72 in39_73 9.241569
Rin39_74 in39_73 in39_74 9.241569
Rin39_75 in39_74 in39_75 9.241569
Rin39_76 in39_75 in39_76 9.241569
Rin39_77 in39_76 in39_77 9.241569
Rin39_78 in39_77 in39_78 9.241569
Rin39_79 in39_78 in39_79 9.241569
Rin39_80 in39_79 in39_80 9.241569
Rin39_81 in39_80 in39_81 9.241569
Rin39_82 in39_81 in39_82 9.241569
Rin39_83 in39_82 in39_83 9.241569
Rin39_84 in39_83 in39_84 9.241569
Rin40_1 in40 in40_1 9.241569
Rin40_2 in40_1 in40_2 9.241569
Rin40_3 in40_2 in40_3 9.241569
Rin40_4 in40_3 in40_4 9.241569
Rin40_5 in40_4 in40_5 9.241569
Rin40_6 in40_5 in40_6 9.241569
Rin40_7 in40_6 in40_7 9.241569
Rin40_8 in40_7 in40_8 9.241569
Rin40_9 in40_8 in40_9 9.241569
Rin40_10 in40_9 in40_10 9.241569
Rin40_11 in40_10 in40_11 9.241569
Rin40_12 in40_11 in40_12 9.241569
Rin40_13 in40_12 in40_13 9.241569
Rin40_14 in40_13 in40_14 9.241569
Rin40_15 in40_14 in40_15 9.241569
Rin40_16 in40_15 in40_16 9.241569
Rin40_17 in40_16 in40_17 9.241569
Rin40_18 in40_17 in40_18 9.241569
Rin40_19 in40_18 in40_19 9.241569
Rin40_20 in40_19 in40_20 9.241569
Rin40_21 in40_20 in40_21 9.241569
Rin40_22 in40_21 in40_22 9.241569
Rin40_23 in40_22 in40_23 9.241569
Rin40_24 in40_23 in40_24 9.241569
Rin40_25 in40_24 in40_25 9.241569
Rin40_26 in40_25 in40_26 9.241569
Rin40_27 in40_26 in40_27 9.241569
Rin40_28 in40_27 in40_28 9.241569
Rin40_29 in40 in40_29 9.241569
Rin40_30 in40_29 in40_30 9.241569
Rin40_31 in40_30 in40_31 9.241569
Rin40_32 in40_31 in40_32 9.241569
Rin40_33 in40_32 in40_33 9.241569
Rin40_34 in40_33 in40_34 9.241569
Rin40_35 in40_34 in40_35 9.241569
Rin40_36 in40_35 in40_36 9.241569
Rin40_37 in40_36 in40_37 9.241569
Rin40_38 in40_37 in40_38 9.241569
Rin40_39 in40_38 in40_39 9.241569
Rin40_40 in40_39 in40_40 9.241569
Rin40_41 in40_40 in40_41 9.241569
Rin40_42 in40_41 in40_42 9.241569
Rin40_43 in40_42 in40_43 9.241569
Rin40_44 in40_43 in40_44 9.241569
Rin40_45 in40_44 in40_45 9.241569
Rin40_46 in40_45 in40_46 9.241569
Rin40_47 in40_46 in40_47 9.241569
Rin40_48 in40_47 in40_48 9.241569
Rin40_49 in40_48 in40_49 9.241569
Rin40_50 in40_49 in40_50 9.241569
Rin40_51 in40_50 in40_51 9.241569
Rin40_52 in40_51 in40_52 9.241569
Rin40_53 in40_52 in40_53 9.241569
Rin40_54 in40_53 in40_54 9.241569
Rin40_55 in40_54 in40_55 9.241569
Rin40_56 in40_55 in40_56 9.241569
Rin40_57 in40 in40_57 9.241569
Rin40_58 in40_57 in40_58 9.241569
Rin40_59 in40_58 in40_59 9.241569
Rin40_60 in40_59 in40_60 9.241569
Rin40_61 in40_60 in40_61 9.241569
Rin40_62 in40_61 in40_62 9.241569
Rin40_63 in40_62 in40_63 9.241569
Rin40_64 in40_63 in40_64 9.241569
Rin40_65 in40_64 in40_65 9.241569
Rin40_66 in40_65 in40_66 9.241569
Rin40_67 in40_66 in40_67 9.241569
Rin40_68 in40_67 in40_68 9.241569
Rin40_69 in40_68 in40_69 9.241569
Rin40_70 in40_69 in40_70 9.241569
Rin40_71 in40_70 in40_71 9.241569
Rin40_72 in40_71 in40_72 9.241569
Rin40_73 in40_72 in40_73 9.241569
Rin40_74 in40_73 in40_74 9.241569
Rin40_75 in40_74 in40_75 9.241569
Rin40_76 in40_75 in40_76 9.241569
Rin40_77 in40_76 in40_77 9.241569
Rin40_78 in40_77 in40_78 9.241569
Rin40_79 in40_78 in40_79 9.241569
Rin40_80 in40_79 in40_80 9.241569
Rin40_81 in40_80 in40_81 9.241569
Rin40_82 in40_81 in40_82 9.241569
Rin40_83 in40_82 in40_83 9.241569
Rin40_84 in40_83 in40_84 9.241569
Rin41_1 in41 in41_1 9.241569
Rin41_2 in41_1 in41_2 9.241569
Rin41_3 in41_2 in41_3 9.241569
Rin41_4 in41_3 in41_4 9.241569
Rin41_5 in41_4 in41_5 9.241569
Rin41_6 in41_5 in41_6 9.241569
Rin41_7 in41_6 in41_7 9.241569
Rin41_8 in41_7 in41_8 9.241569
Rin41_9 in41_8 in41_9 9.241569
Rin41_10 in41_9 in41_10 9.241569
Rin41_11 in41_10 in41_11 9.241569
Rin41_12 in41_11 in41_12 9.241569
Rin41_13 in41_12 in41_13 9.241569
Rin41_14 in41_13 in41_14 9.241569
Rin41_15 in41_14 in41_15 9.241569
Rin41_16 in41_15 in41_16 9.241569
Rin41_17 in41_16 in41_17 9.241569
Rin41_18 in41_17 in41_18 9.241569
Rin41_19 in41_18 in41_19 9.241569
Rin41_20 in41_19 in41_20 9.241569
Rin41_21 in41_20 in41_21 9.241569
Rin41_22 in41_21 in41_22 9.241569
Rin41_23 in41_22 in41_23 9.241569
Rin41_24 in41_23 in41_24 9.241569
Rin41_25 in41_24 in41_25 9.241569
Rin41_26 in41_25 in41_26 9.241569
Rin41_27 in41_26 in41_27 9.241569
Rin41_28 in41_27 in41_28 9.241569
Rin41_29 in41 in41_29 9.241569
Rin41_30 in41_29 in41_30 9.241569
Rin41_31 in41_30 in41_31 9.241569
Rin41_32 in41_31 in41_32 9.241569
Rin41_33 in41_32 in41_33 9.241569
Rin41_34 in41_33 in41_34 9.241569
Rin41_35 in41_34 in41_35 9.241569
Rin41_36 in41_35 in41_36 9.241569
Rin41_37 in41_36 in41_37 9.241569
Rin41_38 in41_37 in41_38 9.241569
Rin41_39 in41_38 in41_39 9.241569
Rin41_40 in41_39 in41_40 9.241569
Rin41_41 in41_40 in41_41 9.241569
Rin41_42 in41_41 in41_42 9.241569
Rin41_43 in41_42 in41_43 9.241569
Rin41_44 in41_43 in41_44 9.241569
Rin41_45 in41_44 in41_45 9.241569
Rin41_46 in41_45 in41_46 9.241569
Rin41_47 in41_46 in41_47 9.241569
Rin41_48 in41_47 in41_48 9.241569
Rin41_49 in41_48 in41_49 9.241569
Rin41_50 in41_49 in41_50 9.241569
Rin41_51 in41_50 in41_51 9.241569
Rin41_52 in41_51 in41_52 9.241569
Rin41_53 in41_52 in41_53 9.241569
Rin41_54 in41_53 in41_54 9.241569
Rin41_55 in41_54 in41_55 9.241569
Rin41_56 in41_55 in41_56 9.241569
Rin41_57 in41 in41_57 9.241569
Rin41_58 in41_57 in41_58 9.241569
Rin41_59 in41_58 in41_59 9.241569
Rin41_60 in41_59 in41_60 9.241569
Rin41_61 in41_60 in41_61 9.241569
Rin41_62 in41_61 in41_62 9.241569
Rin41_63 in41_62 in41_63 9.241569
Rin41_64 in41_63 in41_64 9.241569
Rin41_65 in41_64 in41_65 9.241569
Rin41_66 in41_65 in41_66 9.241569
Rin41_67 in41_66 in41_67 9.241569
Rin41_68 in41_67 in41_68 9.241569
Rin41_69 in41_68 in41_69 9.241569
Rin41_70 in41_69 in41_70 9.241569
Rin41_71 in41_70 in41_71 9.241569
Rin41_72 in41_71 in41_72 9.241569
Rin41_73 in41_72 in41_73 9.241569
Rin41_74 in41_73 in41_74 9.241569
Rin41_75 in41_74 in41_75 9.241569
Rin41_76 in41_75 in41_76 9.241569
Rin41_77 in41_76 in41_77 9.241569
Rin41_78 in41_77 in41_78 9.241569
Rin41_79 in41_78 in41_79 9.241569
Rin41_80 in41_79 in41_80 9.241569
Rin41_81 in41_80 in41_81 9.241569
Rin41_82 in41_81 in41_82 9.241569
Rin41_83 in41_82 in41_83 9.241569
Rin41_84 in41_83 in41_84 9.241569
Rin42_1 in42 in42_1 9.241569
Rin42_2 in42_1 in42_2 9.241569
Rin42_3 in42_2 in42_3 9.241569
Rin42_4 in42_3 in42_4 9.241569
Rin42_5 in42_4 in42_5 9.241569
Rin42_6 in42_5 in42_6 9.241569
Rin42_7 in42_6 in42_7 9.241569
Rin42_8 in42_7 in42_8 9.241569
Rin42_9 in42_8 in42_9 9.241569
Rin42_10 in42_9 in42_10 9.241569
Rin42_11 in42_10 in42_11 9.241569
Rin42_12 in42_11 in42_12 9.241569
Rin42_13 in42_12 in42_13 9.241569
Rin42_14 in42_13 in42_14 9.241569
Rin42_15 in42_14 in42_15 9.241569
Rin42_16 in42_15 in42_16 9.241569
Rin42_17 in42_16 in42_17 9.241569
Rin42_18 in42_17 in42_18 9.241569
Rin42_19 in42_18 in42_19 9.241569
Rin42_20 in42_19 in42_20 9.241569
Rin42_21 in42_20 in42_21 9.241569
Rin42_22 in42_21 in42_22 9.241569
Rin42_23 in42_22 in42_23 9.241569
Rin42_24 in42_23 in42_24 9.241569
Rin42_25 in42_24 in42_25 9.241569
Rin42_26 in42_25 in42_26 9.241569
Rin42_27 in42_26 in42_27 9.241569
Rin42_28 in42_27 in42_28 9.241569
Rin42_29 in42 in42_29 9.241569
Rin42_30 in42_29 in42_30 9.241569
Rin42_31 in42_30 in42_31 9.241569
Rin42_32 in42_31 in42_32 9.241569
Rin42_33 in42_32 in42_33 9.241569
Rin42_34 in42_33 in42_34 9.241569
Rin42_35 in42_34 in42_35 9.241569
Rin42_36 in42_35 in42_36 9.241569
Rin42_37 in42_36 in42_37 9.241569
Rin42_38 in42_37 in42_38 9.241569
Rin42_39 in42_38 in42_39 9.241569
Rin42_40 in42_39 in42_40 9.241569
Rin42_41 in42_40 in42_41 9.241569
Rin42_42 in42_41 in42_42 9.241569
Rin42_43 in42_42 in42_43 9.241569
Rin42_44 in42_43 in42_44 9.241569
Rin42_45 in42_44 in42_45 9.241569
Rin42_46 in42_45 in42_46 9.241569
Rin42_47 in42_46 in42_47 9.241569
Rin42_48 in42_47 in42_48 9.241569
Rin42_49 in42_48 in42_49 9.241569
Rin42_50 in42_49 in42_50 9.241569
Rin42_51 in42_50 in42_51 9.241569
Rin42_52 in42_51 in42_52 9.241569
Rin42_53 in42_52 in42_53 9.241569
Rin42_54 in42_53 in42_54 9.241569
Rin42_55 in42_54 in42_55 9.241569
Rin42_56 in42_55 in42_56 9.241569
Rin42_57 in42 in42_57 9.241569
Rin42_58 in42_57 in42_58 9.241569
Rin42_59 in42_58 in42_59 9.241569
Rin42_60 in42_59 in42_60 9.241569
Rin42_61 in42_60 in42_61 9.241569
Rin42_62 in42_61 in42_62 9.241569
Rin42_63 in42_62 in42_63 9.241569
Rin42_64 in42_63 in42_64 9.241569
Rin42_65 in42_64 in42_65 9.241569
Rin42_66 in42_65 in42_66 9.241569
Rin42_67 in42_66 in42_67 9.241569
Rin42_68 in42_67 in42_68 9.241569
Rin42_69 in42_68 in42_69 9.241569
Rin42_70 in42_69 in42_70 9.241569
Rin42_71 in42_70 in42_71 9.241569
Rin42_72 in42_71 in42_72 9.241569
Rin42_73 in42_72 in42_73 9.241569
Rin42_74 in42_73 in42_74 9.241569
Rin42_75 in42_74 in42_75 9.241569
Rin42_76 in42_75 in42_76 9.241569
Rin42_77 in42_76 in42_77 9.241569
Rin42_78 in42_77 in42_78 9.241569
Rin42_79 in42_78 in42_79 9.241569
Rin42_80 in42_79 in42_80 9.241569
Rin42_81 in42_80 in42_81 9.241569
Rin42_82 in42_81 in42_82 9.241569
Rin42_83 in42_82 in42_83 9.241569
Rin42_84 in42_83 in42_84 9.241569
Rin43_1 in43 in43_1 9.241569
Rin43_2 in43_1 in43_2 9.241569
Rin43_3 in43_2 in43_3 9.241569
Rin43_4 in43_3 in43_4 9.241569
Rin43_5 in43_4 in43_5 9.241569
Rin43_6 in43_5 in43_6 9.241569
Rin43_7 in43_6 in43_7 9.241569
Rin43_8 in43_7 in43_8 9.241569
Rin43_9 in43_8 in43_9 9.241569
Rin43_10 in43_9 in43_10 9.241569
Rin43_11 in43_10 in43_11 9.241569
Rin43_12 in43_11 in43_12 9.241569
Rin43_13 in43_12 in43_13 9.241569
Rin43_14 in43_13 in43_14 9.241569
Rin43_15 in43_14 in43_15 9.241569
Rin43_16 in43_15 in43_16 9.241569
Rin43_17 in43_16 in43_17 9.241569
Rin43_18 in43_17 in43_18 9.241569
Rin43_19 in43_18 in43_19 9.241569
Rin43_20 in43_19 in43_20 9.241569
Rin43_21 in43_20 in43_21 9.241569
Rin43_22 in43_21 in43_22 9.241569
Rin43_23 in43_22 in43_23 9.241569
Rin43_24 in43_23 in43_24 9.241569
Rin43_25 in43_24 in43_25 9.241569
Rin43_26 in43_25 in43_26 9.241569
Rin43_27 in43_26 in43_27 9.241569
Rin43_28 in43_27 in43_28 9.241569
Rin43_29 in43 in43_29 9.241569
Rin43_30 in43_29 in43_30 9.241569
Rin43_31 in43_30 in43_31 9.241569
Rin43_32 in43_31 in43_32 9.241569
Rin43_33 in43_32 in43_33 9.241569
Rin43_34 in43_33 in43_34 9.241569
Rin43_35 in43_34 in43_35 9.241569
Rin43_36 in43_35 in43_36 9.241569
Rin43_37 in43_36 in43_37 9.241569
Rin43_38 in43_37 in43_38 9.241569
Rin43_39 in43_38 in43_39 9.241569
Rin43_40 in43_39 in43_40 9.241569
Rin43_41 in43_40 in43_41 9.241569
Rin43_42 in43_41 in43_42 9.241569
Rin43_43 in43_42 in43_43 9.241569
Rin43_44 in43_43 in43_44 9.241569
Rin43_45 in43_44 in43_45 9.241569
Rin43_46 in43_45 in43_46 9.241569
Rin43_47 in43_46 in43_47 9.241569
Rin43_48 in43_47 in43_48 9.241569
Rin43_49 in43_48 in43_49 9.241569
Rin43_50 in43_49 in43_50 9.241569
Rin43_51 in43_50 in43_51 9.241569
Rin43_52 in43_51 in43_52 9.241569
Rin43_53 in43_52 in43_53 9.241569
Rin43_54 in43_53 in43_54 9.241569
Rin43_55 in43_54 in43_55 9.241569
Rin43_56 in43_55 in43_56 9.241569
Rin43_57 in43 in43_57 9.241569
Rin43_58 in43_57 in43_58 9.241569
Rin43_59 in43_58 in43_59 9.241569
Rin43_60 in43_59 in43_60 9.241569
Rin43_61 in43_60 in43_61 9.241569
Rin43_62 in43_61 in43_62 9.241569
Rin43_63 in43_62 in43_63 9.241569
Rin43_64 in43_63 in43_64 9.241569
Rin43_65 in43_64 in43_65 9.241569
Rin43_66 in43_65 in43_66 9.241569
Rin43_67 in43_66 in43_67 9.241569
Rin43_68 in43_67 in43_68 9.241569
Rin43_69 in43_68 in43_69 9.241569
Rin43_70 in43_69 in43_70 9.241569
Rin43_71 in43_70 in43_71 9.241569
Rin43_72 in43_71 in43_72 9.241569
Rin43_73 in43_72 in43_73 9.241569
Rin43_74 in43_73 in43_74 9.241569
Rin43_75 in43_74 in43_75 9.241569
Rin43_76 in43_75 in43_76 9.241569
Rin43_77 in43_76 in43_77 9.241569
Rin43_78 in43_77 in43_78 9.241569
Rin43_79 in43_78 in43_79 9.241569
Rin43_80 in43_79 in43_80 9.241569
Rin43_81 in43_80 in43_81 9.241569
Rin43_82 in43_81 in43_82 9.241569
Rin43_83 in43_82 in43_83 9.241569
Rin43_84 in43_83 in43_84 9.241569
Rin44_1 in44 in44_1 9.241569
Rin44_2 in44_1 in44_2 9.241569
Rin44_3 in44_2 in44_3 9.241569
Rin44_4 in44_3 in44_4 9.241569
Rin44_5 in44_4 in44_5 9.241569
Rin44_6 in44_5 in44_6 9.241569
Rin44_7 in44_6 in44_7 9.241569
Rin44_8 in44_7 in44_8 9.241569
Rin44_9 in44_8 in44_9 9.241569
Rin44_10 in44_9 in44_10 9.241569
Rin44_11 in44_10 in44_11 9.241569
Rin44_12 in44_11 in44_12 9.241569
Rin44_13 in44_12 in44_13 9.241569
Rin44_14 in44_13 in44_14 9.241569
Rin44_15 in44_14 in44_15 9.241569
Rin44_16 in44_15 in44_16 9.241569
Rin44_17 in44_16 in44_17 9.241569
Rin44_18 in44_17 in44_18 9.241569
Rin44_19 in44_18 in44_19 9.241569
Rin44_20 in44_19 in44_20 9.241569
Rin44_21 in44_20 in44_21 9.241569
Rin44_22 in44_21 in44_22 9.241569
Rin44_23 in44_22 in44_23 9.241569
Rin44_24 in44_23 in44_24 9.241569
Rin44_25 in44_24 in44_25 9.241569
Rin44_26 in44_25 in44_26 9.241569
Rin44_27 in44_26 in44_27 9.241569
Rin44_28 in44_27 in44_28 9.241569
Rin44_29 in44 in44_29 9.241569
Rin44_30 in44_29 in44_30 9.241569
Rin44_31 in44_30 in44_31 9.241569
Rin44_32 in44_31 in44_32 9.241569
Rin44_33 in44_32 in44_33 9.241569
Rin44_34 in44_33 in44_34 9.241569
Rin44_35 in44_34 in44_35 9.241569
Rin44_36 in44_35 in44_36 9.241569
Rin44_37 in44_36 in44_37 9.241569
Rin44_38 in44_37 in44_38 9.241569
Rin44_39 in44_38 in44_39 9.241569
Rin44_40 in44_39 in44_40 9.241569
Rin44_41 in44_40 in44_41 9.241569
Rin44_42 in44_41 in44_42 9.241569
Rin44_43 in44_42 in44_43 9.241569
Rin44_44 in44_43 in44_44 9.241569
Rin44_45 in44_44 in44_45 9.241569
Rin44_46 in44_45 in44_46 9.241569
Rin44_47 in44_46 in44_47 9.241569
Rin44_48 in44_47 in44_48 9.241569
Rin44_49 in44_48 in44_49 9.241569
Rin44_50 in44_49 in44_50 9.241569
Rin44_51 in44_50 in44_51 9.241569
Rin44_52 in44_51 in44_52 9.241569
Rin44_53 in44_52 in44_53 9.241569
Rin44_54 in44_53 in44_54 9.241569
Rin44_55 in44_54 in44_55 9.241569
Rin44_56 in44_55 in44_56 9.241569
Rin44_57 in44 in44_57 9.241569
Rin44_58 in44_57 in44_58 9.241569
Rin44_59 in44_58 in44_59 9.241569
Rin44_60 in44_59 in44_60 9.241569
Rin44_61 in44_60 in44_61 9.241569
Rin44_62 in44_61 in44_62 9.241569
Rin44_63 in44_62 in44_63 9.241569
Rin44_64 in44_63 in44_64 9.241569
Rin44_65 in44_64 in44_65 9.241569
Rin44_66 in44_65 in44_66 9.241569
Rin44_67 in44_66 in44_67 9.241569
Rin44_68 in44_67 in44_68 9.241569
Rin44_69 in44_68 in44_69 9.241569
Rin44_70 in44_69 in44_70 9.241569
Rin44_71 in44_70 in44_71 9.241569
Rin44_72 in44_71 in44_72 9.241569
Rin44_73 in44_72 in44_73 9.241569
Rin44_74 in44_73 in44_74 9.241569
Rin44_75 in44_74 in44_75 9.241569
Rin44_76 in44_75 in44_76 9.241569
Rin44_77 in44_76 in44_77 9.241569
Rin44_78 in44_77 in44_78 9.241569
Rin44_79 in44_78 in44_79 9.241569
Rin44_80 in44_79 in44_80 9.241569
Rin44_81 in44_80 in44_81 9.241569
Rin44_82 in44_81 in44_82 9.241569
Rin44_83 in44_82 in44_83 9.241569
Rin44_84 in44_83 in44_84 9.241569
Rin45_1 in45 in45_1 9.241569
Rin45_2 in45_1 in45_2 9.241569
Rin45_3 in45_2 in45_3 9.241569
Rin45_4 in45_3 in45_4 9.241569
Rin45_5 in45_4 in45_5 9.241569
Rin45_6 in45_5 in45_6 9.241569
Rin45_7 in45_6 in45_7 9.241569
Rin45_8 in45_7 in45_8 9.241569
Rin45_9 in45_8 in45_9 9.241569
Rin45_10 in45_9 in45_10 9.241569
Rin45_11 in45_10 in45_11 9.241569
Rin45_12 in45_11 in45_12 9.241569
Rin45_13 in45_12 in45_13 9.241569
Rin45_14 in45_13 in45_14 9.241569
Rin45_15 in45_14 in45_15 9.241569
Rin45_16 in45_15 in45_16 9.241569
Rin45_17 in45_16 in45_17 9.241569
Rin45_18 in45_17 in45_18 9.241569
Rin45_19 in45_18 in45_19 9.241569
Rin45_20 in45_19 in45_20 9.241569
Rin45_21 in45_20 in45_21 9.241569
Rin45_22 in45_21 in45_22 9.241569
Rin45_23 in45_22 in45_23 9.241569
Rin45_24 in45_23 in45_24 9.241569
Rin45_25 in45_24 in45_25 9.241569
Rin45_26 in45_25 in45_26 9.241569
Rin45_27 in45_26 in45_27 9.241569
Rin45_28 in45_27 in45_28 9.241569
Rin45_29 in45 in45_29 9.241569
Rin45_30 in45_29 in45_30 9.241569
Rin45_31 in45_30 in45_31 9.241569
Rin45_32 in45_31 in45_32 9.241569
Rin45_33 in45_32 in45_33 9.241569
Rin45_34 in45_33 in45_34 9.241569
Rin45_35 in45_34 in45_35 9.241569
Rin45_36 in45_35 in45_36 9.241569
Rin45_37 in45_36 in45_37 9.241569
Rin45_38 in45_37 in45_38 9.241569
Rin45_39 in45_38 in45_39 9.241569
Rin45_40 in45_39 in45_40 9.241569
Rin45_41 in45_40 in45_41 9.241569
Rin45_42 in45_41 in45_42 9.241569
Rin45_43 in45_42 in45_43 9.241569
Rin45_44 in45_43 in45_44 9.241569
Rin45_45 in45_44 in45_45 9.241569
Rin45_46 in45_45 in45_46 9.241569
Rin45_47 in45_46 in45_47 9.241569
Rin45_48 in45_47 in45_48 9.241569
Rin45_49 in45_48 in45_49 9.241569
Rin45_50 in45_49 in45_50 9.241569
Rin45_51 in45_50 in45_51 9.241569
Rin45_52 in45_51 in45_52 9.241569
Rin45_53 in45_52 in45_53 9.241569
Rin45_54 in45_53 in45_54 9.241569
Rin45_55 in45_54 in45_55 9.241569
Rin45_56 in45_55 in45_56 9.241569
Rin45_57 in45 in45_57 9.241569
Rin45_58 in45_57 in45_58 9.241569
Rin45_59 in45_58 in45_59 9.241569
Rin45_60 in45_59 in45_60 9.241569
Rin45_61 in45_60 in45_61 9.241569
Rin45_62 in45_61 in45_62 9.241569
Rin45_63 in45_62 in45_63 9.241569
Rin45_64 in45_63 in45_64 9.241569
Rin45_65 in45_64 in45_65 9.241569
Rin45_66 in45_65 in45_66 9.241569
Rin45_67 in45_66 in45_67 9.241569
Rin45_68 in45_67 in45_68 9.241569
Rin45_69 in45_68 in45_69 9.241569
Rin45_70 in45_69 in45_70 9.241569
Rin45_71 in45_70 in45_71 9.241569
Rin45_72 in45_71 in45_72 9.241569
Rin45_73 in45_72 in45_73 9.241569
Rin45_74 in45_73 in45_74 9.241569
Rin45_75 in45_74 in45_75 9.241569
Rin45_76 in45_75 in45_76 9.241569
Rin45_77 in45_76 in45_77 9.241569
Rin45_78 in45_77 in45_78 9.241569
Rin45_79 in45_78 in45_79 9.241569
Rin45_80 in45_79 in45_80 9.241569
Rin45_81 in45_80 in45_81 9.241569
Rin45_82 in45_81 in45_82 9.241569
Rin45_83 in45_82 in45_83 9.241569
Rin45_84 in45_83 in45_84 9.241569
Rin46_1 in46 in46_1 9.241569
Rin46_2 in46_1 in46_2 9.241569
Rin46_3 in46_2 in46_3 9.241569
Rin46_4 in46_3 in46_4 9.241569
Rin46_5 in46_4 in46_5 9.241569
Rin46_6 in46_5 in46_6 9.241569
Rin46_7 in46_6 in46_7 9.241569
Rin46_8 in46_7 in46_8 9.241569
Rin46_9 in46_8 in46_9 9.241569
Rin46_10 in46_9 in46_10 9.241569
Rin46_11 in46_10 in46_11 9.241569
Rin46_12 in46_11 in46_12 9.241569
Rin46_13 in46_12 in46_13 9.241569
Rin46_14 in46_13 in46_14 9.241569
Rin46_15 in46_14 in46_15 9.241569
Rin46_16 in46_15 in46_16 9.241569
Rin46_17 in46_16 in46_17 9.241569
Rin46_18 in46_17 in46_18 9.241569
Rin46_19 in46_18 in46_19 9.241569
Rin46_20 in46_19 in46_20 9.241569
Rin46_21 in46_20 in46_21 9.241569
Rin46_22 in46_21 in46_22 9.241569
Rin46_23 in46_22 in46_23 9.241569
Rin46_24 in46_23 in46_24 9.241569
Rin46_25 in46_24 in46_25 9.241569
Rin46_26 in46_25 in46_26 9.241569
Rin46_27 in46_26 in46_27 9.241569
Rin46_28 in46_27 in46_28 9.241569
Rin46_29 in46 in46_29 9.241569
Rin46_30 in46_29 in46_30 9.241569
Rin46_31 in46_30 in46_31 9.241569
Rin46_32 in46_31 in46_32 9.241569
Rin46_33 in46_32 in46_33 9.241569
Rin46_34 in46_33 in46_34 9.241569
Rin46_35 in46_34 in46_35 9.241569
Rin46_36 in46_35 in46_36 9.241569
Rin46_37 in46_36 in46_37 9.241569
Rin46_38 in46_37 in46_38 9.241569
Rin46_39 in46_38 in46_39 9.241569
Rin46_40 in46_39 in46_40 9.241569
Rin46_41 in46_40 in46_41 9.241569
Rin46_42 in46_41 in46_42 9.241569
Rin46_43 in46_42 in46_43 9.241569
Rin46_44 in46_43 in46_44 9.241569
Rin46_45 in46_44 in46_45 9.241569
Rin46_46 in46_45 in46_46 9.241569
Rin46_47 in46_46 in46_47 9.241569
Rin46_48 in46_47 in46_48 9.241569
Rin46_49 in46_48 in46_49 9.241569
Rin46_50 in46_49 in46_50 9.241569
Rin46_51 in46_50 in46_51 9.241569
Rin46_52 in46_51 in46_52 9.241569
Rin46_53 in46_52 in46_53 9.241569
Rin46_54 in46_53 in46_54 9.241569
Rin46_55 in46_54 in46_55 9.241569
Rin46_56 in46_55 in46_56 9.241569
Rin46_57 in46 in46_57 9.241569
Rin46_58 in46_57 in46_58 9.241569
Rin46_59 in46_58 in46_59 9.241569
Rin46_60 in46_59 in46_60 9.241569
Rin46_61 in46_60 in46_61 9.241569
Rin46_62 in46_61 in46_62 9.241569
Rin46_63 in46_62 in46_63 9.241569
Rin46_64 in46_63 in46_64 9.241569
Rin46_65 in46_64 in46_65 9.241569
Rin46_66 in46_65 in46_66 9.241569
Rin46_67 in46_66 in46_67 9.241569
Rin46_68 in46_67 in46_68 9.241569
Rin46_69 in46_68 in46_69 9.241569
Rin46_70 in46_69 in46_70 9.241569
Rin46_71 in46_70 in46_71 9.241569
Rin46_72 in46_71 in46_72 9.241569
Rin46_73 in46_72 in46_73 9.241569
Rin46_74 in46_73 in46_74 9.241569
Rin46_75 in46_74 in46_75 9.241569
Rin46_76 in46_75 in46_76 9.241569
Rin46_77 in46_76 in46_77 9.241569
Rin46_78 in46_77 in46_78 9.241569
Rin46_79 in46_78 in46_79 9.241569
Rin46_80 in46_79 in46_80 9.241569
Rin46_81 in46_80 in46_81 9.241569
Rin46_82 in46_81 in46_82 9.241569
Rin46_83 in46_82 in46_83 9.241569
Rin46_84 in46_83 in46_84 9.241569
Rin47_1 in47 in47_1 9.241569
Rin47_2 in47_1 in47_2 9.241569
Rin47_3 in47_2 in47_3 9.241569
Rin47_4 in47_3 in47_4 9.241569
Rin47_5 in47_4 in47_5 9.241569
Rin47_6 in47_5 in47_6 9.241569
Rin47_7 in47_6 in47_7 9.241569
Rin47_8 in47_7 in47_8 9.241569
Rin47_9 in47_8 in47_9 9.241569
Rin47_10 in47_9 in47_10 9.241569
Rin47_11 in47_10 in47_11 9.241569
Rin47_12 in47_11 in47_12 9.241569
Rin47_13 in47_12 in47_13 9.241569
Rin47_14 in47_13 in47_14 9.241569
Rin47_15 in47_14 in47_15 9.241569
Rin47_16 in47_15 in47_16 9.241569
Rin47_17 in47_16 in47_17 9.241569
Rin47_18 in47_17 in47_18 9.241569
Rin47_19 in47_18 in47_19 9.241569
Rin47_20 in47_19 in47_20 9.241569
Rin47_21 in47_20 in47_21 9.241569
Rin47_22 in47_21 in47_22 9.241569
Rin47_23 in47_22 in47_23 9.241569
Rin47_24 in47_23 in47_24 9.241569
Rin47_25 in47_24 in47_25 9.241569
Rin47_26 in47_25 in47_26 9.241569
Rin47_27 in47_26 in47_27 9.241569
Rin47_28 in47_27 in47_28 9.241569
Rin47_29 in47 in47_29 9.241569
Rin47_30 in47_29 in47_30 9.241569
Rin47_31 in47_30 in47_31 9.241569
Rin47_32 in47_31 in47_32 9.241569
Rin47_33 in47_32 in47_33 9.241569
Rin47_34 in47_33 in47_34 9.241569
Rin47_35 in47_34 in47_35 9.241569
Rin47_36 in47_35 in47_36 9.241569
Rin47_37 in47_36 in47_37 9.241569
Rin47_38 in47_37 in47_38 9.241569
Rin47_39 in47_38 in47_39 9.241569
Rin47_40 in47_39 in47_40 9.241569
Rin47_41 in47_40 in47_41 9.241569
Rin47_42 in47_41 in47_42 9.241569
Rin47_43 in47_42 in47_43 9.241569
Rin47_44 in47_43 in47_44 9.241569
Rin47_45 in47_44 in47_45 9.241569
Rin47_46 in47_45 in47_46 9.241569
Rin47_47 in47_46 in47_47 9.241569
Rin47_48 in47_47 in47_48 9.241569
Rin47_49 in47_48 in47_49 9.241569
Rin47_50 in47_49 in47_50 9.241569
Rin47_51 in47_50 in47_51 9.241569
Rin47_52 in47_51 in47_52 9.241569
Rin47_53 in47_52 in47_53 9.241569
Rin47_54 in47_53 in47_54 9.241569
Rin47_55 in47_54 in47_55 9.241569
Rin47_56 in47_55 in47_56 9.241569
Rin47_57 in47 in47_57 9.241569
Rin47_58 in47_57 in47_58 9.241569
Rin47_59 in47_58 in47_59 9.241569
Rin47_60 in47_59 in47_60 9.241569
Rin47_61 in47_60 in47_61 9.241569
Rin47_62 in47_61 in47_62 9.241569
Rin47_63 in47_62 in47_63 9.241569
Rin47_64 in47_63 in47_64 9.241569
Rin47_65 in47_64 in47_65 9.241569
Rin47_66 in47_65 in47_66 9.241569
Rin47_67 in47_66 in47_67 9.241569
Rin47_68 in47_67 in47_68 9.241569
Rin47_69 in47_68 in47_69 9.241569
Rin47_70 in47_69 in47_70 9.241569
Rin47_71 in47_70 in47_71 9.241569
Rin47_72 in47_71 in47_72 9.241569
Rin47_73 in47_72 in47_73 9.241569
Rin47_74 in47_73 in47_74 9.241569
Rin47_75 in47_74 in47_75 9.241569
Rin47_76 in47_75 in47_76 9.241569
Rin47_77 in47_76 in47_77 9.241569
Rin47_78 in47_77 in47_78 9.241569
Rin47_79 in47_78 in47_79 9.241569
Rin47_80 in47_79 in47_80 9.241569
Rin47_81 in47_80 in47_81 9.241569
Rin47_82 in47_81 in47_82 9.241569
Rin47_83 in47_82 in47_83 9.241569
Rin47_84 in47_83 in47_84 9.241569
Rin48_1 in48 in48_1 9.241569
Rin48_2 in48_1 in48_2 9.241569
Rin48_3 in48_2 in48_3 9.241569
Rin48_4 in48_3 in48_4 9.241569
Rin48_5 in48_4 in48_5 9.241569
Rin48_6 in48_5 in48_6 9.241569
Rin48_7 in48_6 in48_7 9.241569
Rin48_8 in48_7 in48_8 9.241569
Rin48_9 in48_8 in48_9 9.241569
Rin48_10 in48_9 in48_10 9.241569
Rin48_11 in48_10 in48_11 9.241569
Rin48_12 in48_11 in48_12 9.241569
Rin48_13 in48_12 in48_13 9.241569
Rin48_14 in48_13 in48_14 9.241569
Rin48_15 in48_14 in48_15 9.241569
Rin48_16 in48_15 in48_16 9.241569
Rin48_17 in48_16 in48_17 9.241569
Rin48_18 in48_17 in48_18 9.241569
Rin48_19 in48_18 in48_19 9.241569
Rin48_20 in48_19 in48_20 9.241569
Rin48_21 in48_20 in48_21 9.241569
Rin48_22 in48_21 in48_22 9.241569
Rin48_23 in48_22 in48_23 9.241569
Rin48_24 in48_23 in48_24 9.241569
Rin48_25 in48_24 in48_25 9.241569
Rin48_26 in48_25 in48_26 9.241569
Rin48_27 in48_26 in48_27 9.241569
Rin48_28 in48_27 in48_28 9.241569
Rin48_29 in48 in48_29 9.241569
Rin48_30 in48_29 in48_30 9.241569
Rin48_31 in48_30 in48_31 9.241569
Rin48_32 in48_31 in48_32 9.241569
Rin48_33 in48_32 in48_33 9.241569
Rin48_34 in48_33 in48_34 9.241569
Rin48_35 in48_34 in48_35 9.241569
Rin48_36 in48_35 in48_36 9.241569
Rin48_37 in48_36 in48_37 9.241569
Rin48_38 in48_37 in48_38 9.241569
Rin48_39 in48_38 in48_39 9.241569
Rin48_40 in48_39 in48_40 9.241569
Rin48_41 in48_40 in48_41 9.241569
Rin48_42 in48_41 in48_42 9.241569
Rin48_43 in48_42 in48_43 9.241569
Rin48_44 in48_43 in48_44 9.241569
Rin48_45 in48_44 in48_45 9.241569
Rin48_46 in48_45 in48_46 9.241569
Rin48_47 in48_46 in48_47 9.241569
Rin48_48 in48_47 in48_48 9.241569
Rin48_49 in48_48 in48_49 9.241569
Rin48_50 in48_49 in48_50 9.241569
Rin48_51 in48_50 in48_51 9.241569
Rin48_52 in48_51 in48_52 9.241569
Rin48_53 in48_52 in48_53 9.241569
Rin48_54 in48_53 in48_54 9.241569
Rin48_55 in48_54 in48_55 9.241569
Rin48_56 in48_55 in48_56 9.241569
Rin48_57 in48 in48_57 9.241569
Rin48_58 in48_57 in48_58 9.241569
Rin48_59 in48_58 in48_59 9.241569
Rin48_60 in48_59 in48_60 9.241569
Rin48_61 in48_60 in48_61 9.241569
Rin48_62 in48_61 in48_62 9.241569
Rin48_63 in48_62 in48_63 9.241569
Rin48_64 in48_63 in48_64 9.241569
Rin48_65 in48_64 in48_65 9.241569
Rin48_66 in48_65 in48_66 9.241569
Rin48_67 in48_66 in48_67 9.241569
Rin48_68 in48_67 in48_68 9.241569
Rin48_69 in48_68 in48_69 9.241569
Rin48_70 in48_69 in48_70 9.241569
Rin48_71 in48_70 in48_71 9.241569
Rin48_72 in48_71 in48_72 9.241569
Rin48_73 in48_72 in48_73 9.241569
Rin48_74 in48_73 in48_74 9.241569
Rin48_75 in48_74 in48_75 9.241569
Rin48_76 in48_75 in48_76 9.241569
Rin48_77 in48_76 in48_77 9.241569
Rin48_78 in48_77 in48_78 9.241569
Rin48_79 in48_78 in48_79 9.241569
Rin48_80 in48_79 in48_80 9.241569
Rin48_81 in48_80 in48_81 9.241569
Rin48_82 in48_81 in48_82 9.241569
Rin48_83 in48_82 in48_83 9.241569
Rin48_84 in48_83 in48_84 9.241569
Rin49_1 in49 in49_1 9.241569
Rin49_2 in49_1 in49_2 9.241569
Rin49_3 in49_2 in49_3 9.241569
Rin49_4 in49_3 in49_4 9.241569
Rin49_5 in49_4 in49_5 9.241569
Rin49_6 in49_5 in49_6 9.241569
Rin49_7 in49_6 in49_7 9.241569
Rin49_8 in49_7 in49_8 9.241569
Rin49_9 in49_8 in49_9 9.241569
Rin49_10 in49_9 in49_10 9.241569
Rin49_11 in49_10 in49_11 9.241569
Rin49_12 in49_11 in49_12 9.241569
Rin49_13 in49_12 in49_13 9.241569
Rin49_14 in49_13 in49_14 9.241569
Rin49_15 in49_14 in49_15 9.241569
Rin49_16 in49_15 in49_16 9.241569
Rin49_17 in49_16 in49_17 9.241569
Rin49_18 in49_17 in49_18 9.241569
Rin49_19 in49_18 in49_19 9.241569
Rin49_20 in49_19 in49_20 9.241569
Rin49_21 in49_20 in49_21 9.241569
Rin49_22 in49_21 in49_22 9.241569
Rin49_23 in49_22 in49_23 9.241569
Rin49_24 in49_23 in49_24 9.241569
Rin49_25 in49_24 in49_25 9.241569
Rin49_26 in49_25 in49_26 9.241569
Rin49_27 in49_26 in49_27 9.241569
Rin49_28 in49_27 in49_28 9.241569
Rin49_29 in49 in49_29 9.241569
Rin49_30 in49_29 in49_30 9.241569
Rin49_31 in49_30 in49_31 9.241569
Rin49_32 in49_31 in49_32 9.241569
Rin49_33 in49_32 in49_33 9.241569
Rin49_34 in49_33 in49_34 9.241569
Rin49_35 in49_34 in49_35 9.241569
Rin49_36 in49_35 in49_36 9.241569
Rin49_37 in49_36 in49_37 9.241569
Rin49_38 in49_37 in49_38 9.241569
Rin49_39 in49_38 in49_39 9.241569
Rin49_40 in49_39 in49_40 9.241569
Rin49_41 in49_40 in49_41 9.241569
Rin49_42 in49_41 in49_42 9.241569
Rin49_43 in49_42 in49_43 9.241569
Rin49_44 in49_43 in49_44 9.241569
Rin49_45 in49_44 in49_45 9.241569
Rin49_46 in49_45 in49_46 9.241569
Rin49_47 in49_46 in49_47 9.241569
Rin49_48 in49_47 in49_48 9.241569
Rin49_49 in49_48 in49_49 9.241569
Rin49_50 in49_49 in49_50 9.241569
Rin49_51 in49_50 in49_51 9.241569
Rin49_52 in49_51 in49_52 9.241569
Rin49_53 in49_52 in49_53 9.241569
Rin49_54 in49_53 in49_54 9.241569
Rin49_55 in49_54 in49_55 9.241569
Rin49_56 in49_55 in49_56 9.241569
Rin49_57 in49 in49_57 9.241569
Rin49_58 in49_57 in49_58 9.241569
Rin49_59 in49_58 in49_59 9.241569
Rin49_60 in49_59 in49_60 9.241569
Rin49_61 in49_60 in49_61 9.241569
Rin49_62 in49_61 in49_62 9.241569
Rin49_63 in49_62 in49_63 9.241569
Rin49_64 in49_63 in49_64 9.241569
Rin49_65 in49_64 in49_65 9.241569
Rin49_66 in49_65 in49_66 9.241569
Rin49_67 in49_66 in49_67 9.241569
Rin49_68 in49_67 in49_68 9.241569
Rin49_69 in49_68 in49_69 9.241569
Rin49_70 in49_69 in49_70 9.241569
Rin49_71 in49_70 in49_71 9.241569
Rin49_72 in49_71 in49_72 9.241569
Rin49_73 in49_72 in49_73 9.241569
Rin49_74 in49_73 in49_74 9.241569
Rin49_75 in49_74 in49_75 9.241569
Rin49_76 in49_75 in49_76 9.241569
Rin49_77 in49_76 in49_77 9.241569
Rin49_78 in49_77 in49_78 9.241569
Rin49_79 in49_78 in49_79 9.241569
Rin49_80 in49_79 in49_80 9.241569
Rin49_81 in49_80 in49_81 9.241569
Rin49_82 in49_81 in49_82 9.241569
Rin49_83 in49_82 in49_83 9.241569
Rin49_84 in49_83 in49_84 9.241569
Rin50_1 in50 in50_1 9.241569
Rin50_2 in50_1 in50_2 9.241569
Rin50_3 in50_2 in50_3 9.241569
Rin50_4 in50_3 in50_4 9.241569
Rin50_5 in50_4 in50_5 9.241569
Rin50_6 in50_5 in50_6 9.241569
Rin50_7 in50_6 in50_7 9.241569
Rin50_8 in50_7 in50_8 9.241569
Rin50_9 in50_8 in50_9 9.241569
Rin50_10 in50_9 in50_10 9.241569
Rin50_11 in50_10 in50_11 9.241569
Rin50_12 in50_11 in50_12 9.241569
Rin50_13 in50_12 in50_13 9.241569
Rin50_14 in50_13 in50_14 9.241569
Rin50_15 in50_14 in50_15 9.241569
Rin50_16 in50_15 in50_16 9.241569
Rin50_17 in50_16 in50_17 9.241569
Rin50_18 in50_17 in50_18 9.241569
Rin50_19 in50_18 in50_19 9.241569
Rin50_20 in50_19 in50_20 9.241569
Rin50_21 in50_20 in50_21 9.241569
Rin50_22 in50_21 in50_22 9.241569
Rin50_23 in50_22 in50_23 9.241569
Rin50_24 in50_23 in50_24 9.241569
Rin50_25 in50_24 in50_25 9.241569
Rin50_26 in50_25 in50_26 9.241569
Rin50_27 in50_26 in50_27 9.241569
Rin50_28 in50_27 in50_28 9.241569
Rin50_29 in50 in50_29 9.241569
Rin50_30 in50_29 in50_30 9.241569
Rin50_31 in50_30 in50_31 9.241569
Rin50_32 in50_31 in50_32 9.241569
Rin50_33 in50_32 in50_33 9.241569
Rin50_34 in50_33 in50_34 9.241569
Rin50_35 in50_34 in50_35 9.241569
Rin50_36 in50_35 in50_36 9.241569
Rin50_37 in50_36 in50_37 9.241569
Rin50_38 in50_37 in50_38 9.241569
Rin50_39 in50_38 in50_39 9.241569
Rin50_40 in50_39 in50_40 9.241569
Rin50_41 in50_40 in50_41 9.241569
Rin50_42 in50_41 in50_42 9.241569
Rin50_43 in50_42 in50_43 9.241569
Rin50_44 in50_43 in50_44 9.241569
Rin50_45 in50_44 in50_45 9.241569
Rin50_46 in50_45 in50_46 9.241569
Rin50_47 in50_46 in50_47 9.241569
Rin50_48 in50_47 in50_48 9.241569
Rin50_49 in50_48 in50_49 9.241569
Rin50_50 in50_49 in50_50 9.241569
Rin50_51 in50_50 in50_51 9.241569
Rin50_52 in50_51 in50_52 9.241569
Rin50_53 in50_52 in50_53 9.241569
Rin50_54 in50_53 in50_54 9.241569
Rin50_55 in50_54 in50_55 9.241569
Rin50_56 in50_55 in50_56 9.241569
Rin50_57 in50 in50_57 9.241569
Rin50_58 in50_57 in50_58 9.241569
Rin50_59 in50_58 in50_59 9.241569
Rin50_60 in50_59 in50_60 9.241569
Rin50_61 in50_60 in50_61 9.241569
Rin50_62 in50_61 in50_62 9.241569
Rin50_63 in50_62 in50_63 9.241569
Rin50_64 in50_63 in50_64 9.241569
Rin50_65 in50_64 in50_65 9.241569
Rin50_66 in50_65 in50_66 9.241569
Rin50_67 in50_66 in50_67 9.241569
Rin50_68 in50_67 in50_68 9.241569
Rin50_69 in50_68 in50_69 9.241569
Rin50_70 in50_69 in50_70 9.241569
Rin50_71 in50_70 in50_71 9.241569
Rin50_72 in50_71 in50_72 9.241569
Rin50_73 in50_72 in50_73 9.241569
Rin50_74 in50_73 in50_74 9.241569
Rin50_75 in50_74 in50_75 9.241569
Rin50_76 in50_75 in50_76 9.241569
Rin50_77 in50_76 in50_77 9.241569
Rin50_78 in50_77 in50_78 9.241569
Rin50_79 in50_78 in50_79 9.241569
Rin50_80 in50_79 in50_80 9.241569
Rin50_81 in50_80 in50_81 9.241569
Rin50_82 in50_81 in50_82 9.241569
Rin50_83 in50_82 in50_83 9.241569
Rin50_84 in50_83 in50_84 9.241569
Rin51_1 in51 in51_1 9.241569
Rin51_2 in51_1 in51_2 9.241569
Rin51_3 in51_2 in51_3 9.241569
Rin51_4 in51_3 in51_4 9.241569
Rin51_5 in51_4 in51_5 9.241569
Rin51_6 in51_5 in51_6 9.241569
Rin51_7 in51_6 in51_7 9.241569
Rin51_8 in51_7 in51_8 9.241569
Rin51_9 in51_8 in51_9 9.241569
Rin51_10 in51_9 in51_10 9.241569
Rin51_11 in51_10 in51_11 9.241569
Rin51_12 in51_11 in51_12 9.241569
Rin51_13 in51_12 in51_13 9.241569
Rin51_14 in51_13 in51_14 9.241569
Rin51_15 in51_14 in51_15 9.241569
Rin51_16 in51_15 in51_16 9.241569
Rin51_17 in51_16 in51_17 9.241569
Rin51_18 in51_17 in51_18 9.241569
Rin51_19 in51_18 in51_19 9.241569
Rin51_20 in51_19 in51_20 9.241569
Rin51_21 in51_20 in51_21 9.241569
Rin51_22 in51_21 in51_22 9.241569
Rin51_23 in51_22 in51_23 9.241569
Rin51_24 in51_23 in51_24 9.241569
Rin51_25 in51_24 in51_25 9.241569
Rin51_26 in51_25 in51_26 9.241569
Rin51_27 in51_26 in51_27 9.241569
Rin51_28 in51_27 in51_28 9.241569
Rin51_29 in51 in51_29 9.241569
Rin51_30 in51_29 in51_30 9.241569
Rin51_31 in51_30 in51_31 9.241569
Rin51_32 in51_31 in51_32 9.241569
Rin51_33 in51_32 in51_33 9.241569
Rin51_34 in51_33 in51_34 9.241569
Rin51_35 in51_34 in51_35 9.241569
Rin51_36 in51_35 in51_36 9.241569
Rin51_37 in51_36 in51_37 9.241569
Rin51_38 in51_37 in51_38 9.241569
Rin51_39 in51_38 in51_39 9.241569
Rin51_40 in51_39 in51_40 9.241569
Rin51_41 in51_40 in51_41 9.241569
Rin51_42 in51_41 in51_42 9.241569
Rin51_43 in51_42 in51_43 9.241569
Rin51_44 in51_43 in51_44 9.241569
Rin51_45 in51_44 in51_45 9.241569
Rin51_46 in51_45 in51_46 9.241569
Rin51_47 in51_46 in51_47 9.241569
Rin51_48 in51_47 in51_48 9.241569
Rin51_49 in51_48 in51_49 9.241569
Rin51_50 in51_49 in51_50 9.241569
Rin51_51 in51_50 in51_51 9.241569
Rin51_52 in51_51 in51_52 9.241569
Rin51_53 in51_52 in51_53 9.241569
Rin51_54 in51_53 in51_54 9.241569
Rin51_55 in51_54 in51_55 9.241569
Rin51_56 in51_55 in51_56 9.241569
Rin51_57 in51 in51_57 9.241569
Rin51_58 in51_57 in51_58 9.241569
Rin51_59 in51_58 in51_59 9.241569
Rin51_60 in51_59 in51_60 9.241569
Rin51_61 in51_60 in51_61 9.241569
Rin51_62 in51_61 in51_62 9.241569
Rin51_63 in51_62 in51_63 9.241569
Rin51_64 in51_63 in51_64 9.241569
Rin51_65 in51_64 in51_65 9.241569
Rin51_66 in51_65 in51_66 9.241569
Rin51_67 in51_66 in51_67 9.241569
Rin51_68 in51_67 in51_68 9.241569
Rin51_69 in51_68 in51_69 9.241569
Rin51_70 in51_69 in51_70 9.241569
Rin51_71 in51_70 in51_71 9.241569
Rin51_72 in51_71 in51_72 9.241569
Rin51_73 in51_72 in51_73 9.241569
Rin51_74 in51_73 in51_74 9.241569
Rin51_75 in51_74 in51_75 9.241569
Rin51_76 in51_75 in51_76 9.241569
Rin51_77 in51_76 in51_77 9.241569
Rin51_78 in51_77 in51_78 9.241569
Rin51_79 in51_78 in51_79 9.241569
Rin51_80 in51_79 in51_80 9.241569
Rin51_81 in51_80 in51_81 9.241569
Rin51_82 in51_81 in51_82 9.241569
Rin51_83 in51_82 in51_83 9.241569
Rin51_84 in51_83 in51_84 9.241569
Rin52_1 in52 in52_1 9.241569
Rin52_2 in52_1 in52_2 9.241569
Rin52_3 in52_2 in52_3 9.241569
Rin52_4 in52_3 in52_4 9.241569
Rin52_5 in52_4 in52_5 9.241569
Rin52_6 in52_5 in52_6 9.241569
Rin52_7 in52_6 in52_7 9.241569
Rin52_8 in52_7 in52_8 9.241569
Rin52_9 in52_8 in52_9 9.241569
Rin52_10 in52_9 in52_10 9.241569
Rin52_11 in52_10 in52_11 9.241569
Rin52_12 in52_11 in52_12 9.241569
Rin52_13 in52_12 in52_13 9.241569
Rin52_14 in52_13 in52_14 9.241569
Rin52_15 in52_14 in52_15 9.241569
Rin52_16 in52_15 in52_16 9.241569
Rin52_17 in52_16 in52_17 9.241569
Rin52_18 in52_17 in52_18 9.241569
Rin52_19 in52_18 in52_19 9.241569
Rin52_20 in52_19 in52_20 9.241569
Rin52_21 in52_20 in52_21 9.241569
Rin52_22 in52_21 in52_22 9.241569
Rin52_23 in52_22 in52_23 9.241569
Rin52_24 in52_23 in52_24 9.241569
Rin52_25 in52_24 in52_25 9.241569
Rin52_26 in52_25 in52_26 9.241569
Rin52_27 in52_26 in52_27 9.241569
Rin52_28 in52_27 in52_28 9.241569
Rin52_29 in52 in52_29 9.241569
Rin52_30 in52_29 in52_30 9.241569
Rin52_31 in52_30 in52_31 9.241569
Rin52_32 in52_31 in52_32 9.241569
Rin52_33 in52_32 in52_33 9.241569
Rin52_34 in52_33 in52_34 9.241569
Rin52_35 in52_34 in52_35 9.241569
Rin52_36 in52_35 in52_36 9.241569
Rin52_37 in52_36 in52_37 9.241569
Rin52_38 in52_37 in52_38 9.241569
Rin52_39 in52_38 in52_39 9.241569
Rin52_40 in52_39 in52_40 9.241569
Rin52_41 in52_40 in52_41 9.241569
Rin52_42 in52_41 in52_42 9.241569
Rin52_43 in52_42 in52_43 9.241569
Rin52_44 in52_43 in52_44 9.241569
Rin52_45 in52_44 in52_45 9.241569
Rin52_46 in52_45 in52_46 9.241569
Rin52_47 in52_46 in52_47 9.241569
Rin52_48 in52_47 in52_48 9.241569
Rin52_49 in52_48 in52_49 9.241569
Rin52_50 in52_49 in52_50 9.241569
Rin52_51 in52_50 in52_51 9.241569
Rin52_52 in52_51 in52_52 9.241569
Rin52_53 in52_52 in52_53 9.241569
Rin52_54 in52_53 in52_54 9.241569
Rin52_55 in52_54 in52_55 9.241569
Rin52_56 in52_55 in52_56 9.241569
Rin52_57 in52 in52_57 9.241569
Rin52_58 in52_57 in52_58 9.241569
Rin52_59 in52_58 in52_59 9.241569
Rin52_60 in52_59 in52_60 9.241569
Rin52_61 in52_60 in52_61 9.241569
Rin52_62 in52_61 in52_62 9.241569
Rin52_63 in52_62 in52_63 9.241569
Rin52_64 in52_63 in52_64 9.241569
Rin52_65 in52_64 in52_65 9.241569
Rin52_66 in52_65 in52_66 9.241569
Rin52_67 in52_66 in52_67 9.241569
Rin52_68 in52_67 in52_68 9.241569
Rin52_69 in52_68 in52_69 9.241569
Rin52_70 in52_69 in52_70 9.241569
Rin52_71 in52_70 in52_71 9.241569
Rin52_72 in52_71 in52_72 9.241569
Rin52_73 in52_72 in52_73 9.241569
Rin52_74 in52_73 in52_74 9.241569
Rin52_75 in52_74 in52_75 9.241569
Rin52_76 in52_75 in52_76 9.241569
Rin52_77 in52_76 in52_77 9.241569
Rin52_78 in52_77 in52_78 9.241569
Rin52_79 in52_78 in52_79 9.241569
Rin52_80 in52_79 in52_80 9.241569
Rin52_81 in52_80 in52_81 9.241569
Rin52_82 in52_81 in52_82 9.241569
Rin52_83 in52_82 in52_83 9.241569
Rin52_84 in52_83 in52_84 9.241569
Rin53_1 in53 in53_1 9.241569
Rin53_2 in53_1 in53_2 9.241569
Rin53_3 in53_2 in53_3 9.241569
Rin53_4 in53_3 in53_4 9.241569
Rin53_5 in53_4 in53_5 9.241569
Rin53_6 in53_5 in53_6 9.241569
Rin53_7 in53_6 in53_7 9.241569
Rin53_8 in53_7 in53_8 9.241569
Rin53_9 in53_8 in53_9 9.241569
Rin53_10 in53_9 in53_10 9.241569
Rin53_11 in53_10 in53_11 9.241569
Rin53_12 in53_11 in53_12 9.241569
Rin53_13 in53_12 in53_13 9.241569
Rin53_14 in53_13 in53_14 9.241569
Rin53_15 in53_14 in53_15 9.241569
Rin53_16 in53_15 in53_16 9.241569
Rin53_17 in53_16 in53_17 9.241569
Rin53_18 in53_17 in53_18 9.241569
Rin53_19 in53_18 in53_19 9.241569
Rin53_20 in53_19 in53_20 9.241569
Rin53_21 in53_20 in53_21 9.241569
Rin53_22 in53_21 in53_22 9.241569
Rin53_23 in53_22 in53_23 9.241569
Rin53_24 in53_23 in53_24 9.241569
Rin53_25 in53_24 in53_25 9.241569
Rin53_26 in53_25 in53_26 9.241569
Rin53_27 in53_26 in53_27 9.241569
Rin53_28 in53_27 in53_28 9.241569
Rin53_29 in53 in53_29 9.241569
Rin53_30 in53_29 in53_30 9.241569
Rin53_31 in53_30 in53_31 9.241569
Rin53_32 in53_31 in53_32 9.241569
Rin53_33 in53_32 in53_33 9.241569
Rin53_34 in53_33 in53_34 9.241569
Rin53_35 in53_34 in53_35 9.241569
Rin53_36 in53_35 in53_36 9.241569
Rin53_37 in53_36 in53_37 9.241569
Rin53_38 in53_37 in53_38 9.241569
Rin53_39 in53_38 in53_39 9.241569
Rin53_40 in53_39 in53_40 9.241569
Rin53_41 in53_40 in53_41 9.241569
Rin53_42 in53_41 in53_42 9.241569
Rin53_43 in53_42 in53_43 9.241569
Rin53_44 in53_43 in53_44 9.241569
Rin53_45 in53_44 in53_45 9.241569
Rin53_46 in53_45 in53_46 9.241569
Rin53_47 in53_46 in53_47 9.241569
Rin53_48 in53_47 in53_48 9.241569
Rin53_49 in53_48 in53_49 9.241569
Rin53_50 in53_49 in53_50 9.241569
Rin53_51 in53_50 in53_51 9.241569
Rin53_52 in53_51 in53_52 9.241569
Rin53_53 in53_52 in53_53 9.241569
Rin53_54 in53_53 in53_54 9.241569
Rin53_55 in53_54 in53_55 9.241569
Rin53_56 in53_55 in53_56 9.241569
Rin53_57 in53 in53_57 9.241569
Rin53_58 in53_57 in53_58 9.241569
Rin53_59 in53_58 in53_59 9.241569
Rin53_60 in53_59 in53_60 9.241569
Rin53_61 in53_60 in53_61 9.241569
Rin53_62 in53_61 in53_62 9.241569
Rin53_63 in53_62 in53_63 9.241569
Rin53_64 in53_63 in53_64 9.241569
Rin53_65 in53_64 in53_65 9.241569
Rin53_66 in53_65 in53_66 9.241569
Rin53_67 in53_66 in53_67 9.241569
Rin53_68 in53_67 in53_68 9.241569
Rin53_69 in53_68 in53_69 9.241569
Rin53_70 in53_69 in53_70 9.241569
Rin53_71 in53_70 in53_71 9.241569
Rin53_72 in53_71 in53_72 9.241569
Rin53_73 in53_72 in53_73 9.241569
Rin53_74 in53_73 in53_74 9.241569
Rin53_75 in53_74 in53_75 9.241569
Rin53_76 in53_75 in53_76 9.241569
Rin53_77 in53_76 in53_77 9.241569
Rin53_78 in53_77 in53_78 9.241569
Rin53_79 in53_78 in53_79 9.241569
Rin53_80 in53_79 in53_80 9.241569
Rin53_81 in53_80 in53_81 9.241569
Rin53_82 in53_81 in53_82 9.241569
Rin53_83 in53_82 in53_83 9.241569
Rin53_84 in53_83 in53_84 9.241569
Rin54_1 in54 in54_1 9.241569
Rin54_2 in54_1 in54_2 9.241569
Rin54_3 in54_2 in54_3 9.241569
Rin54_4 in54_3 in54_4 9.241569
Rin54_5 in54_4 in54_5 9.241569
Rin54_6 in54_5 in54_6 9.241569
Rin54_7 in54_6 in54_7 9.241569
Rin54_8 in54_7 in54_8 9.241569
Rin54_9 in54_8 in54_9 9.241569
Rin54_10 in54_9 in54_10 9.241569
Rin54_11 in54_10 in54_11 9.241569
Rin54_12 in54_11 in54_12 9.241569
Rin54_13 in54_12 in54_13 9.241569
Rin54_14 in54_13 in54_14 9.241569
Rin54_15 in54_14 in54_15 9.241569
Rin54_16 in54_15 in54_16 9.241569
Rin54_17 in54_16 in54_17 9.241569
Rin54_18 in54_17 in54_18 9.241569
Rin54_19 in54_18 in54_19 9.241569
Rin54_20 in54_19 in54_20 9.241569
Rin54_21 in54_20 in54_21 9.241569
Rin54_22 in54_21 in54_22 9.241569
Rin54_23 in54_22 in54_23 9.241569
Rin54_24 in54_23 in54_24 9.241569
Rin54_25 in54_24 in54_25 9.241569
Rin54_26 in54_25 in54_26 9.241569
Rin54_27 in54_26 in54_27 9.241569
Rin54_28 in54_27 in54_28 9.241569
Rin54_29 in54 in54_29 9.241569
Rin54_30 in54_29 in54_30 9.241569
Rin54_31 in54_30 in54_31 9.241569
Rin54_32 in54_31 in54_32 9.241569
Rin54_33 in54_32 in54_33 9.241569
Rin54_34 in54_33 in54_34 9.241569
Rin54_35 in54_34 in54_35 9.241569
Rin54_36 in54_35 in54_36 9.241569
Rin54_37 in54_36 in54_37 9.241569
Rin54_38 in54_37 in54_38 9.241569
Rin54_39 in54_38 in54_39 9.241569
Rin54_40 in54_39 in54_40 9.241569
Rin54_41 in54_40 in54_41 9.241569
Rin54_42 in54_41 in54_42 9.241569
Rin54_43 in54_42 in54_43 9.241569
Rin54_44 in54_43 in54_44 9.241569
Rin54_45 in54_44 in54_45 9.241569
Rin54_46 in54_45 in54_46 9.241569
Rin54_47 in54_46 in54_47 9.241569
Rin54_48 in54_47 in54_48 9.241569
Rin54_49 in54_48 in54_49 9.241569
Rin54_50 in54_49 in54_50 9.241569
Rin54_51 in54_50 in54_51 9.241569
Rin54_52 in54_51 in54_52 9.241569
Rin54_53 in54_52 in54_53 9.241569
Rin54_54 in54_53 in54_54 9.241569
Rin54_55 in54_54 in54_55 9.241569
Rin54_56 in54_55 in54_56 9.241569
Rin54_57 in54 in54_57 9.241569
Rin54_58 in54_57 in54_58 9.241569
Rin54_59 in54_58 in54_59 9.241569
Rin54_60 in54_59 in54_60 9.241569
Rin54_61 in54_60 in54_61 9.241569
Rin54_62 in54_61 in54_62 9.241569
Rin54_63 in54_62 in54_63 9.241569
Rin54_64 in54_63 in54_64 9.241569
Rin54_65 in54_64 in54_65 9.241569
Rin54_66 in54_65 in54_66 9.241569
Rin54_67 in54_66 in54_67 9.241569
Rin54_68 in54_67 in54_68 9.241569
Rin54_69 in54_68 in54_69 9.241569
Rin54_70 in54_69 in54_70 9.241569
Rin54_71 in54_70 in54_71 9.241569
Rin54_72 in54_71 in54_72 9.241569
Rin54_73 in54_72 in54_73 9.241569
Rin54_74 in54_73 in54_74 9.241569
Rin54_75 in54_74 in54_75 9.241569
Rin54_76 in54_75 in54_76 9.241569
Rin54_77 in54_76 in54_77 9.241569
Rin54_78 in54_77 in54_78 9.241569
Rin54_79 in54_78 in54_79 9.241569
Rin54_80 in54_79 in54_80 9.241569
Rin54_81 in54_80 in54_81 9.241569
Rin54_82 in54_81 in54_82 9.241569
Rin54_83 in54_82 in54_83 9.241569
Rin54_84 in54_83 in54_84 9.241569
Rin55_1 in55 in55_1 9.241569
Rin55_2 in55_1 in55_2 9.241569
Rin55_3 in55_2 in55_3 9.241569
Rin55_4 in55_3 in55_4 9.241569
Rin55_5 in55_4 in55_5 9.241569
Rin55_6 in55_5 in55_6 9.241569
Rin55_7 in55_6 in55_7 9.241569
Rin55_8 in55_7 in55_8 9.241569
Rin55_9 in55_8 in55_9 9.241569
Rin55_10 in55_9 in55_10 9.241569
Rin55_11 in55_10 in55_11 9.241569
Rin55_12 in55_11 in55_12 9.241569
Rin55_13 in55_12 in55_13 9.241569
Rin55_14 in55_13 in55_14 9.241569
Rin55_15 in55_14 in55_15 9.241569
Rin55_16 in55_15 in55_16 9.241569
Rin55_17 in55_16 in55_17 9.241569
Rin55_18 in55_17 in55_18 9.241569
Rin55_19 in55_18 in55_19 9.241569
Rin55_20 in55_19 in55_20 9.241569
Rin55_21 in55_20 in55_21 9.241569
Rin55_22 in55_21 in55_22 9.241569
Rin55_23 in55_22 in55_23 9.241569
Rin55_24 in55_23 in55_24 9.241569
Rin55_25 in55_24 in55_25 9.241569
Rin55_26 in55_25 in55_26 9.241569
Rin55_27 in55_26 in55_27 9.241569
Rin55_28 in55_27 in55_28 9.241569
Rin55_29 in55 in55_29 9.241569
Rin55_30 in55_29 in55_30 9.241569
Rin55_31 in55_30 in55_31 9.241569
Rin55_32 in55_31 in55_32 9.241569
Rin55_33 in55_32 in55_33 9.241569
Rin55_34 in55_33 in55_34 9.241569
Rin55_35 in55_34 in55_35 9.241569
Rin55_36 in55_35 in55_36 9.241569
Rin55_37 in55_36 in55_37 9.241569
Rin55_38 in55_37 in55_38 9.241569
Rin55_39 in55_38 in55_39 9.241569
Rin55_40 in55_39 in55_40 9.241569
Rin55_41 in55_40 in55_41 9.241569
Rin55_42 in55_41 in55_42 9.241569
Rin55_43 in55_42 in55_43 9.241569
Rin55_44 in55_43 in55_44 9.241569
Rin55_45 in55_44 in55_45 9.241569
Rin55_46 in55_45 in55_46 9.241569
Rin55_47 in55_46 in55_47 9.241569
Rin55_48 in55_47 in55_48 9.241569
Rin55_49 in55_48 in55_49 9.241569
Rin55_50 in55_49 in55_50 9.241569
Rin55_51 in55_50 in55_51 9.241569
Rin55_52 in55_51 in55_52 9.241569
Rin55_53 in55_52 in55_53 9.241569
Rin55_54 in55_53 in55_54 9.241569
Rin55_55 in55_54 in55_55 9.241569
Rin55_56 in55_55 in55_56 9.241569
Rin55_57 in55 in55_57 9.241569
Rin55_58 in55_57 in55_58 9.241569
Rin55_59 in55_58 in55_59 9.241569
Rin55_60 in55_59 in55_60 9.241569
Rin55_61 in55_60 in55_61 9.241569
Rin55_62 in55_61 in55_62 9.241569
Rin55_63 in55_62 in55_63 9.241569
Rin55_64 in55_63 in55_64 9.241569
Rin55_65 in55_64 in55_65 9.241569
Rin55_66 in55_65 in55_66 9.241569
Rin55_67 in55_66 in55_67 9.241569
Rin55_68 in55_67 in55_68 9.241569
Rin55_69 in55_68 in55_69 9.241569
Rin55_70 in55_69 in55_70 9.241569
Rin55_71 in55_70 in55_71 9.241569
Rin55_72 in55_71 in55_72 9.241569
Rin55_73 in55_72 in55_73 9.241569
Rin55_74 in55_73 in55_74 9.241569
Rin55_75 in55_74 in55_75 9.241569
Rin55_76 in55_75 in55_76 9.241569
Rin55_77 in55_76 in55_77 9.241569
Rin55_78 in55_77 in55_78 9.241569
Rin55_79 in55_78 in55_79 9.241569
Rin55_80 in55_79 in55_80 9.241569
Rin55_81 in55_80 in55_81 9.241569
Rin55_82 in55_81 in55_82 9.241569
Rin55_83 in55_82 in55_83 9.241569
Rin55_84 in55_83 in55_84 9.241569
Rin56_1 in56 in56_1 9.241569
Rin56_2 in56_1 in56_2 9.241569
Rin56_3 in56_2 in56_3 9.241569
Rin56_4 in56_3 in56_4 9.241569
Rin56_5 in56_4 in56_5 9.241569
Rin56_6 in56_5 in56_6 9.241569
Rin56_7 in56_6 in56_7 9.241569
Rin56_8 in56_7 in56_8 9.241569
Rin56_9 in56_8 in56_9 9.241569
Rin56_10 in56_9 in56_10 9.241569
Rin56_11 in56_10 in56_11 9.241569
Rin56_12 in56_11 in56_12 9.241569
Rin56_13 in56_12 in56_13 9.241569
Rin56_14 in56_13 in56_14 9.241569
Rin56_15 in56_14 in56_15 9.241569
Rin56_16 in56_15 in56_16 9.241569
Rin56_17 in56_16 in56_17 9.241569
Rin56_18 in56_17 in56_18 9.241569
Rin56_19 in56_18 in56_19 9.241569
Rin56_20 in56_19 in56_20 9.241569
Rin56_21 in56_20 in56_21 9.241569
Rin56_22 in56_21 in56_22 9.241569
Rin56_23 in56_22 in56_23 9.241569
Rin56_24 in56_23 in56_24 9.241569
Rin56_25 in56_24 in56_25 9.241569
Rin56_26 in56_25 in56_26 9.241569
Rin56_27 in56_26 in56_27 9.241569
Rin56_28 in56_27 in56_28 9.241569
Rin56_29 in56 in56_29 9.241569
Rin56_30 in56_29 in56_30 9.241569
Rin56_31 in56_30 in56_31 9.241569
Rin56_32 in56_31 in56_32 9.241569
Rin56_33 in56_32 in56_33 9.241569
Rin56_34 in56_33 in56_34 9.241569
Rin56_35 in56_34 in56_35 9.241569
Rin56_36 in56_35 in56_36 9.241569
Rin56_37 in56_36 in56_37 9.241569
Rin56_38 in56_37 in56_38 9.241569
Rin56_39 in56_38 in56_39 9.241569
Rin56_40 in56_39 in56_40 9.241569
Rin56_41 in56_40 in56_41 9.241569
Rin56_42 in56_41 in56_42 9.241569
Rin56_43 in56_42 in56_43 9.241569
Rin56_44 in56_43 in56_44 9.241569
Rin56_45 in56_44 in56_45 9.241569
Rin56_46 in56_45 in56_46 9.241569
Rin56_47 in56_46 in56_47 9.241569
Rin56_48 in56_47 in56_48 9.241569
Rin56_49 in56_48 in56_49 9.241569
Rin56_50 in56_49 in56_50 9.241569
Rin56_51 in56_50 in56_51 9.241569
Rin56_52 in56_51 in56_52 9.241569
Rin56_53 in56_52 in56_53 9.241569
Rin56_54 in56_53 in56_54 9.241569
Rin56_55 in56_54 in56_55 9.241569
Rin56_56 in56_55 in56_56 9.241569
Rin56_57 in56 in56_57 9.241569
Rin56_58 in56_57 in56_58 9.241569
Rin56_59 in56_58 in56_59 9.241569
Rin56_60 in56_59 in56_60 9.241569
Rin56_61 in56_60 in56_61 9.241569
Rin56_62 in56_61 in56_62 9.241569
Rin56_63 in56_62 in56_63 9.241569
Rin56_64 in56_63 in56_64 9.241569
Rin56_65 in56_64 in56_65 9.241569
Rin56_66 in56_65 in56_66 9.241569
Rin56_67 in56_66 in56_67 9.241569
Rin56_68 in56_67 in56_68 9.241569
Rin56_69 in56_68 in56_69 9.241569
Rin56_70 in56_69 in56_70 9.241569
Rin56_71 in56_70 in56_71 9.241569
Rin56_72 in56_71 in56_72 9.241569
Rin56_73 in56_72 in56_73 9.241569
Rin56_74 in56_73 in56_74 9.241569
Rin56_75 in56_74 in56_75 9.241569
Rin56_76 in56_75 in56_76 9.241569
Rin56_77 in56_76 in56_77 9.241569
Rin56_78 in56_77 in56_78 9.241569
Rin56_79 in56_78 in56_79 9.241569
Rin56_80 in56_79 in56_80 9.241569
Rin56_81 in56_80 in56_81 9.241569
Rin56_82 in56_81 in56_82 9.241569
Rin56_83 in56_82 in56_83 9.241569
Rin56_84 in56_83 in56_84 9.241569
Rin57_1 in57 in57_1 9.241569
Rin57_2 in57_1 in57_2 9.241569
Rin57_3 in57_2 in57_3 9.241569
Rin57_4 in57_3 in57_4 9.241569
Rin57_5 in57_4 in57_5 9.241569
Rin57_6 in57_5 in57_6 9.241569
Rin57_7 in57_6 in57_7 9.241569
Rin57_8 in57_7 in57_8 9.241569
Rin57_9 in57_8 in57_9 9.241569
Rin57_10 in57_9 in57_10 9.241569
Rin57_11 in57_10 in57_11 9.241569
Rin57_12 in57_11 in57_12 9.241569
Rin57_13 in57_12 in57_13 9.241569
Rin57_14 in57_13 in57_14 9.241569
Rin57_15 in57_14 in57_15 9.241569
Rin57_16 in57_15 in57_16 9.241569
Rin57_17 in57_16 in57_17 9.241569
Rin57_18 in57_17 in57_18 9.241569
Rin57_19 in57_18 in57_19 9.241569
Rin57_20 in57_19 in57_20 9.241569
Rin57_21 in57_20 in57_21 9.241569
Rin57_22 in57_21 in57_22 9.241569
Rin57_23 in57_22 in57_23 9.241569
Rin57_24 in57_23 in57_24 9.241569
Rin57_25 in57_24 in57_25 9.241569
Rin57_26 in57_25 in57_26 9.241569
Rin57_27 in57_26 in57_27 9.241569
Rin57_28 in57_27 in57_28 9.241569
Rin57_29 in57 in57_29 9.241569
Rin57_30 in57_29 in57_30 9.241569
Rin57_31 in57_30 in57_31 9.241569
Rin57_32 in57_31 in57_32 9.241569
Rin57_33 in57_32 in57_33 9.241569
Rin57_34 in57_33 in57_34 9.241569
Rin57_35 in57_34 in57_35 9.241569
Rin57_36 in57_35 in57_36 9.241569
Rin57_37 in57_36 in57_37 9.241569
Rin57_38 in57_37 in57_38 9.241569
Rin57_39 in57_38 in57_39 9.241569
Rin57_40 in57_39 in57_40 9.241569
Rin57_41 in57_40 in57_41 9.241569
Rin57_42 in57_41 in57_42 9.241569
Rin57_43 in57_42 in57_43 9.241569
Rin57_44 in57_43 in57_44 9.241569
Rin57_45 in57_44 in57_45 9.241569
Rin57_46 in57_45 in57_46 9.241569
Rin57_47 in57_46 in57_47 9.241569
Rin57_48 in57_47 in57_48 9.241569
Rin57_49 in57_48 in57_49 9.241569
Rin57_50 in57_49 in57_50 9.241569
Rin57_51 in57_50 in57_51 9.241569
Rin57_52 in57_51 in57_52 9.241569
Rin57_53 in57_52 in57_53 9.241569
Rin57_54 in57_53 in57_54 9.241569
Rin57_55 in57_54 in57_55 9.241569
Rin57_56 in57_55 in57_56 9.241569
Rin57_57 in57 in57_57 9.241569
Rin57_58 in57_57 in57_58 9.241569
Rin57_59 in57_58 in57_59 9.241569
Rin57_60 in57_59 in57_60 9.241569
Rin57_61 in57_60 in57_61 9.241569
Rin57_62 in57_61 in57_62 9.241569
Rin57_63 in57_62 in57_63 9.241569
Rin57_64 in57_63 in57_64 9.241569
Rin57_65 in57_64 in57_65 9.241569
Rin57_66 in57_65 in57_66 9.241569
Rin57_67 in57_66 in57_67 9.241569
Rin57_68 in57_67 in57_68 9.241569
Rin57_69 in57_68 in57_69 9.241569
Rin57_70 in57_69 in57_70 9.241569
Rin57_71 in57_70 in57_71 9.241569
Rin57_72 in57_71 in57_72 9.241569
Rin57_73 in57_72 in57_73 9.241569
Rin57_74 in57_73 in57_74 9.241569
Rin57_75 in57_74 in57_75 9.241569
Rin57_76 in57_75 in57_76 9.241569
Rin57_77 in57_76 in57_77 9.241569
Rin57_78 in57_77 in57_78 9.241569
Rin57_79 in57_78 in57_79 9.241569
Rin57_80 in57_79 in57_80 9.241569
Rin57_81 in57_80 in57_81 9.241569
Rin57_82 in57_81 in57_82 9.241569
Rin57_83 in57_82 in57_83 9.241569
Rin57_84 in57_83 in57_84 9.241569
Rin58_1 in58 in58_1 9.241569
Rin58_2 in58_1 in58_2 9.241569
Rin58_3 in58_2 in58_3 9.241569
Rin58_4 in58_3 in58_4 9.241569
Rin58_5 in58_4 in58_5 9.241569
Rin58_6 in58_5 in58_6 9.241569
Rin58_7 in58_6 in58_7 9.241569
Rin58_8 in58_7 in58_8 9.241569
Rin58_9 in58_8 in58_9 9.241569
Rin58_10 in58_9 in58_10 9.241569
Rin58_11 in58_10 in58_11 9.241569
Rin58_12 in58_11 in58_12 9.241569
Rin58_13 in58_12 in58_13 9.241569
Rin58_14 in58_13 in58_14 9.241569
Rin58_15 in58_14 in58_15 9.241569
Rin58_16 in58_15 in58_16 9.241569
Rin58_17 in58_16 in58_17 9.241569
Rin58_18 in58_17 in58_18 9.241569
Rin58_19 in58_18 in58_19 9.241569
Rin58_20 in58_19 in58_20 9.241569
Rin58_21 in58_20 in58_21 9.241569
Rin58_22 in58_21 in58_22 9.241569
Rin58_23 in58_22 in58_23 9.241569
Rin58_24 in58_23 in58_24 9.241569
Rin58_25 in58_24 in58_25 9.241569
Rin58_26 in58_25 in58_26 9.241569
Rin58_27 in58_26 in58_27 9.241569
Rin58_28 in58_27 in58_28 9.241569
Rin58_29 in58 in58_29 9.241569
Rin58_30 in58_29 in58_30 9.241569
Rin58_31 in58_30 in58_31 9.241569
Rin58_32 in58_31 in58_32 9.241569
Rin58_33 in58_32 in58_33 9.241569
Rin58_34 in58_33 in58_34 9.241569
Rin58_35 in58_34 in58_35 9.241569
Rin58_36 in58_35 in58_36 9.241569
Rin58_37 in58_36 in58_37 9.241569
Rin58_38 in58_37 in58_38 9.241569
Rin58_39 in58_38 in58_39 9.241569
Rin58_40 in58_39 in58_40 9.241569
Rin58_41 in58_40 in58_41 9.241569
Rin58_42 in58_41 in58_42 9.241569
Rin58_43 in58_42 in58_43 9.241569
Rin58_44 in58_43 in58_44 9.241569
Rin58_45 in58_44 in58_45 9.241569
Rin58_46 in58_45 in58_46 9.241569
Rin58_47 in58_46 in58_47 9.241569
Rin58_48 in58_47 in58_48 9.241569
Rin58_49 in58_48 in58_49 9.241569
Rin58_50 in58_49 in58_50 9.241569
Rin58_51 in58_50 in58_51 9.241569
Rin58_52 in58_51 in58_52 9.241569
Rin58_53 in58_52 in58_53 9.241569
Rin58_54 in58_53 in58_54 9.241569
Rin58_55 in58_54 in58_55 9.241569
Rin58_56 in58_55 in58_56 9.241569
Rin58_57 in58 in58_57 9.241569
Rin58_58 in58_57 in58_58 9.241569
Rin58_59 in58_58 in58_59 9.241569
Rin58_60 in58_59 in58_60 9.241569
Rin58_61 in58_60 in58_61 9.241569
Rin58_62 in58_61 in58_62 9.241569
Rin58_63 in58_62 in58_63 9.241569
Rin58_64 in58_63 in58_64 9.241569
Rin58_65 in58_64 in58_65 9.241569
Rin58_66 in58_65 in58_66 9.241569
Rin58_67 in58_66 in58_67 9.241569
Rin58_68 in58_67 in58_68 9.241569
Rin58_69 in58_68 in58_69 9.241569
Rin58_70 in58_69 in58_70 9.241569
Rin58_71 in58_70 in58_71 9.241569
Rin58_72 in58_71 in58_72 9.241569
Rin58_73 in58_72 in58_73 9.241569
Rin58_74 in58_73 in58_74 9.241569
Rin58_75 in58_74 in58_75 9.241569
Rin58_76 in58_75 in58_76 9.241569
Rin58_77 in58_76 in58_77 9.241569
Rin58_78 in58_77 in58_78 9.241569
Rin58_79 in58_78 in58_79 9.241569
Rin58_80 in58_79 in58_80 9.241569
Rin58_81 in58_80 in58_81 9.241569
Rin58_82 in58_81 in58_82 9.241569
Rin58_83 in58_82 in58_83 9.241569
Rin58_84 in58_83 in58_84 9.241569
Rin59_1 in59 in59_1 9.241569
Rin59_2 in59_1 in59_2 9.241569
Rin59_3 in59_2 in59_3 9.241569
Rin59_4 in59_3 in59_4 9.241569
Rin59_5 in59_4 in59_5 9.241569
Rin59_6 in59_5 in59_6 9.241569
Rin59_7 in59_6 in59_7 9.241569
Rin59_8 in59_7 in59_8 9.241569
Rin59_9 in59_8 in59_9 9.241569
Rin59_10 in59_9 in59_10 9.241569
Rin59_11 in59_10 in59_11 9.241569
Rin59_12 in59_11 in59_12 9.241569
Rin59_13 in59_12 in59_13 9.241569
Rin59_14 in59_13 in59_14 9.241569
Rin59_15 in59_14 in59_15 9.241569
Rin59_16 in59_15 in59_16 9.241569
Rin59_17 in59_16 in59_17 9.241569
Rin59_18 in59_17 in59_18 9.241569
Rin59_19 in59_18 in59_19 9.241569
Rin59_20 in59_19 in59_20 9.241569
Rin59_21 in59_20 in59_21 9.241569
Rin59_22 in59_21 in59_22 9.241569
Rin59_23 in59_22 in59_23 9.241569
Rin59_24 in59_23 in59_24 9.241569
Rin59_25 in59_24 in59_25 9.241569
Rin59_26 in59_25 in59_26 9.241569
Rin59_27 in59_26 in59_27 9.241569
Rin59_28 in59_27 in59_28 9.241569
Rin59_29 in59 in59_29 9.241569
Rin59_30 in59_29 in59_30 9.241569
Rin59_31 in59_30 in59_31 9.241569
Rin59_32 in59_31 in59_32 9.241569
Rin59_33 in59_32 in59_33 9.241569
Rin59_34 in59_33 in59_34 9.241569
Rin59_35 in59_34 in59_35 9.241569
Rin59_36 in59_35 in59_36 9.241569
Rin59_37 in59_36 in59_37 9.241569
Rin59_38 in59_37 in59_38 9.241569
Rin59_39 in59_38 in59_39 9.241569
Rin59_40 in59_39 in59_40 9.241569
Rin59_41 in59_40 in59_41 9.241569
Rin59_42 in59_41 in59_42 9.241569
Rin59_43 in59_42 in59_43 9.241569
Rin59_44 in59_43 in59_44 9.241569
Rin59_45 in59_44 in59_45 9.241569
Rin59_46 in59_45 in59_46 9.241569
Rin59_47 in59_46 in59_47 9.241569
Rin59_48 in59_47 in59_48 9.241569
Rin59_49 in59_48 in59_49 9.241569
Rin59_50 in59_49 in59_50 9.241569
Rin59_51 in59_50 in59_51 9.241569
Rin59_52 in59_51 in59_52 9.241569
Rin59_53 in59_52 in59_53 9.241569
Rin59_54 in59_53 in59_54 9.241569
Rin59_55 in59_54 in59_55 9.241569
Rin59_56 in59_55 in59_56 9.241569
Rin59_57 in59 in59_57 9.241569
Rin59_58 in59_57 in59_58 9.241569
Rin59_59 in59_58 in59_59 9.241569
Rin59_60 in59_59 in59_60 9.241569
Rin59_61 in59_60 in59_61 9.241569
Rin59_62 in59_61 in59_62 9.241569
Rin59_63 in59_62 in59_63 9.241569
Rin59_64 in59_63 in59_64 9.241569
Rin59_65 in59_64 in59_65 9.241569
Rin59_66 in59_65 in59_66 9.241569
Rin59_67 in59_66 in59_67 9.241569
Rin59_68 in59_67 in59_68 9.241569
Rin59_69 in59_68 in59_69 9.241569
Rin59_70 in59_69 in59_70 9.241569
Rin59_71 in59_70 in59_71 9.241569
Rin59_72 in59_71 in59_72 9.241569
Rin59_73 in59_72 in59_73 9.241569
Rin59_74 in59_73 in59_74 9.241569
Rin59_75 in59_74 in59_75 9.241569
Rin59_76 in59_75 in59_76 9.241569
Rin59_77 in59_76 in59_77 9.241569
Rin59_78 in59_77 in59_78 9.241569
Rin59_79 in59_78 in59_79 9.241569
Rin59_80 in59_79 in59_80 9.241569
Rin59_81 in59_80 in59_81 9.241569
Rin59_82 in59_81 in59_82 9.241569
Rin59_83 in59_82 in59_83 9.241569
Rin59_84 in59_83 in59_84 9.241569
Rin60_1 in60 in60_1 9.241569
Rin60_2 in60_1 in60_2 9.241569
Rin60_3 in60_2 in60_3 9.241569
Rin60_4 in60_3 in60_4 9.241569
Rin60_5 in60_4 in60_5 9.241569
Rin60_6 in60_5 in60_6 9.241569
Rin60_7 in60_6 in60_7 9.241569
Rin60_8 in60_7 in60_8 9.241569
Rin60_9 in60_8 in60_9 9.241569
Rin60_10 in60_9 in60_10 9.241569
Rin60_11 in60_10 in60_11 9.241569
Rin60_12 in60_11 in60_12 9.241569
Rin60_13 in60_12 in60_13 9.241569
Rin60_14 in60_13 in60_14 9.241569
Rin60_15 in60_14 in60_15 9.241569
Rin60_16 in60_15 in60_16 9.241569
Rin60_17 in60_16 in60_17 9.241569
Rin60_18 in60_17 in60_18 9.241569
Rin60_19 in60_18 in60_19 9.241569
Rin60_20 in60_19 in60_20 9.241569
Rin60_21 in60_20 in60_21 9.241569
Rin60_22 in60_21 in60_22 9.241569
Rin60_23 in60_22 in60_23 9.241569
Rin60_24 in60_23 in60_24 9.241569
Rin60_25 in60_24 in60_25 9.241569
Rin60_26 in60_25 in60_26 9.241569
Rin60_27 in60_26 in60_27 9.241569
Rin60_28 in60_27 in60_28 9.241569
Rin60_29 in60 in60_29 9.241569
Rin60_30 in60_29 in60_30 9.241569
Rin60_31 in60_30 in60_31 9.241569
Rin60_32 in60_31 in60_32 9.241569
Rin60_33 in60_32 in60_33 9.241569
Rin60_34 in60_33 in60_34 9.241569
Rin60_35 in60_34 in60_35 9.241569
Rin60_36 in60_35 in60_36 9.241569
Rin60_37 in60_36 in60_37 9.241569
Rin60_38 in60_37 in60_38 9.241569
Rin60_39 in60_38 in60_39 9.241569
Rin60_40 in60_39 in60_40 9.241569
Rin60_41 in60_40 in60_41 9.241569
Rin60_42 in60_41 in60_42 9.241569
Rin60_43 in60_42 in60_43 9.241569
Rin60_44 in60_43 in60_44 9.241569
Rin60_45 in60_44 in60_45 9.241569
Rin60_46 in60_45 in60_46 9.241569
Rin60_47 in60_46 in60_47 9.241569
Rin60_48 in60_47 in60_48 9.241569
Rin60_49 in60_48 in60_49 9.241569
Rin60_50 in60_49 in60_50 9.241569
Rin60_51 in60_50 in60_51 9.241569
Rin60_52 in60_51 in60_52 9.241569
Rin60_53 in60_52 in60_53 9.241569
Rin60_54 in60_53 in60_54 9.241569
Rin60_55 in60_54 in60_55 9.241569
Rin60_56 in60_55 in60_56 9.241569
Rin60_57 in60 in60_57 9.241569
Rin60_58 in60_57 in60_58 9.241569
Rin60_59 in60_58 in60_59 9.241569
Rin60_60 in60_59 in60_60 9.241569
Rin60_61 in60_60 in60_61 9.241569
Rin60_62 in60_61 in60_62 9.241569
Rin60_63 in60_62 in60_63 9.241569
Rin60_64 in60_63 in60_64 9.241569
Rin60_65 in60_64 in60_65 9.241569
Rin60_66 in60_65 in60_66 9.241569
Rin60_67 in60_66 in60_67 9.241569
Rin60_68 in60_67 in60_68 9.241569
Rin60_69 in60_68 in60_69 9.241569
Rin60_70 in60_69 in60_70 9.241569
Rin60_71 in60_70 in60_71 9.241569
Rin60_72 in60_71 in60_72 9.241569
Rin60_73 in60_72 in60_73 9.241569
Rin60_74 in60_73 in60_74 9.241569
Rin60_75 in60_74 in60_75 9.241569
Rin60_76 in60_75 in60_76 9.241569
Rin60_77 in60_76 in60_77 9.241569
Rin60_78 in60_77 in60_78 9.241569
Rin60_79 in60_78 in60_79 9.241569
Rin60_80 in60_79 in60_80 9.241569
Rin60_81 in60_80 in60_81 9.241569
Rin60_82 in60_81 in60_82 9.241569
Rin60_83 in60_82 in60_83 9.241569
Rin60_84 in60_83 in60_84 9.241569
Rin61_1 in61 in61_1 9.241569
Rin61_2 in61_1 in61_2 9.241569
Rin61_3 in61_2 in61_3 9.241569
Rin61_4 in61_3 in61_4 9.241569
Rin61_5 in61_4 in61_5 9.241569
Rin61_6 in61_5 in61_6 9.241569
Rin61_7 in61_6 in61_7 9.241569
Rin61_8 in61_7 in61_8 9.241569
Rin61_9 in61_8 in61_9 9.241569
Rin61_10 in61_9 in61_10 9.241569
Rin61_11 in61_10 in61_11 9.241569
Rin61_12 in61_11 in61_12 9.241569
Rin61_13 in61_12 in61_13 9.241569
Rin61_14 in61_13 in61_14 9.241569
Rin61_15 in61_14 in61_15 9.241569
Rin61_16 in61_15 in61_16 9.241569
Rin61_17 in61_16 in61_17 9.241569
Rin61_18 in61_17 in61_18 9.241569
Rin61_19 in61_18 in61_19 9.241569
Rin61_20 in61_19 in61_20 9.241569
Rin61_21 in61_20 in61_21 9.241569
Rin61_22 in61_21 in61_22 9.241569
Rin61_23 in61_22 in61_23 9.241569
Rin61_24 in61_23 in61_24 9.241569
Rin61_25 in61_24 in61_25 9.241569
Rin61_26 in61_25 in61_26 9.241569
Rin61_27 in61_26 in61_27 9.241569
Rin61_28 in61_27 in61_28 9.241569
Rin61_29 in61 in61_29 9.241569
Rin61_30 in61_29 in61_30 9.241569
Rin61_31 in61_30 in61_31 9.241569
Rin61_32 in61_31 in61_32 9.241569
Rin61_33 in61_32 in61_33 9.241569
Rin61_34 in61_33 in61_34 9.241569
Rin61_35 in61_34 in61_35 9.241569
Rin61_36 in61_35 in61_36 9.241569
Rin61_37 in61_36 in61_37 9.241569
Rin61_38 in61_37 in61_38 9.241569
Rin61_39 in61_38 in61_39 9.241569
Rin61_40 in61_39 in61_40 9.241569
Rin61_41 in61_40 in61_41 9.241569
Rin61_42 in61_41 in61_42 9.241569
Rin61_43 in61_42 in61_43 9.241569
Rin61_44 in61_43 in61_44 9.241569
Rin61_45 in61_44 in61_45 9.241569
Rin61_46 in61_45 in61_46 9.241569
Rin61_47 in61_46 in61_47 9.241569
Rin61_48 in61_47 in61_48 9.241569
Rin61_49 in61_48 in61_49 9.241569
Rin61_50 in61_49 in61_50 9.241569
Rin61_51 in61_50 in61_51 9.241569
Rin61_52 in61_51 in61_52 9.241569
Rin61_53 in61_52 in61_53 9.241569
Rin61_54 in61_53 in61_54 9.241569
Rin61_55 in61_54 in61_55 9.241569
Rin61_56 in61_55 in61_56 9.241569
Rin61_57 in61 in61_57 9.241569
Rin61_58 in61_57 in61_58 9.241569
Rin61_59 in61_58 in61_59 9.241569
Rin61_60 in61_59 in61_60 9.241569
Rin61_61 in61_60 in61_61 9.241569
Rin61_62 in61_61 in61_62 9.241569
Rin61_63 in61_62 in61_63 9.241569
Rin61_64 in61_63 in61_64 9.241569
Rin61_65 in61_64 in61_65 9.241569
Rin61_66 in61_65 in61_66 9.241569
Rin61_67 in61_66 in61_67 9.241569
Rin61_68 in61_67 in61_68 9.241569
Rin61_69 in61_68 in61_69 9.241569
Rin61_70 in61_69 in61_70 9.241569
Rin61_71 in61_70 in61_71 9.241569
Rin61_72 in61_71 in61_72 9.241569
Rin61_73 in61_72 in61_73 9.241569
Rin61_74 in61_73 in61_74 9.241569
Rin61_75 in61_74 in61_75 9.241569
Rin61_76 in61_75 in61_76 9.241569
Rin61_77 in61_76 in61_77 9.241569
Rin61_78 in61_77 in61_78 9.241569
Rin61_79 in61_78 in61_79 9.241569
Rin61_80 in61_79 in61_80 9.241569
Rin61_81 in61_80 in61_81 9.241569
Rin61_82 in61_81 in61_82 9.241569
Rin61_83 in61_82 in61_83 9.241569
Rin61_84 in61_83 in61_84 9.241569
Rin62_1 in62 in62_1 9.241569
Rin62_2 in62_1 in62_2 9.241569
Rin62_3 in62_2 in62_3 9.241569
Rin62_4 in62_3 in62_4 9.241569
Rin62_5 in62_4 in62_5 9.241569
Rin62_6 in62_5 in62_6 9.241569
Rin62_7 in62_6 in62_7 9.241569
Rin62_8 in62_7 in62_8 9.241569
Rin62_9 in62_8 in62_9 9.241569
Rin62_10 in62_9 in62_10 9.241569
Rin62_11 in62_10 in62_11 9.241569
Rin62_12 in62_11 in62_12 9.241569
Rin62_13 in62_12 in62_13 9.241569
Rin62_14 in62_13 in62_14 9.241569
Rin62_15 in62_14 in62_15 9.241569
Rin62_16 in62_15 in62_16 9.241569
Rin62_17 in62_16 in62_17 9.241569
Rin62_18 in62_17 in62_18 9.241569
Rin62_19 in62_18 in62_19 9.241569
Rin62_20 in62_19 in62_20 9.241569
Rin62_21 in62_20 in62_21 9.241569
Rin62_22 in62_21 in62_22 9.241569
Rin62_23 in62_22 in62_23 9.241569
Rin62_24 in62_23 in62_24 9.241569
Rin62_25 in62_24 in62_25 9.241569
Rin62_26 in62_25 in62_26 9.241569
Rin62_27 in62_26 in62_27 9.241569
Rin62_28 in62_27 in62_28 9.241569
Rin62_29 in62 in62_29 9.241569
Rin62_30 in62_29 in62_30 9.241569
Rin62_31 in62_30 in62_31 9.241569
Rin62_32 in62_31 in62_32 9.241569
Rin62_33 in62_32 in62_33 9.241569
Rin62_34 in62_33 in62_34 9.241569
Rin62_35 in62_34 in62_35 9.241569
Rin62_36 in62_35 in62_36 9.241569
Rin62_37 in62_36 in62_37 9.241569
Rin62_38 in62_37 in62_38 9.241569
Rin62_39 in62_38 in62_39 9.241569
Rin62_40 in62_39 in62_40 9.241569
Rin62_41 in62_40 in62_41 9.241569
Rin62_42 in62_41 in62_42 9.241569
Rin62_43 in62_42 in62_43 9.241569
Rin62_44 in62_43 in62_44 9.241569
Rin62_45 in62_44 in62_45 9.241569
Rin62_46 in62_45 in62_46 9.241569
Rin62_47 in62_46 in62_47 9.241569
Rin62_48 in62_47 in62_48 9.241569
Rin62_49 in62_48 in62_49 9.241569
Rin62_50 in62_49 in62_50 9.241569
Rin62_51 in62_50 in62_51 9.241569
Rin62_52 in62_51 in62_52 9.241569
Rin62_53 in62_52 in62_53 9.241569
Rin62_54 in62_53 in62_54 9.241569
Rin62_55 in62_54 in62_55 9.241569
Rin62_56 in62_55 in62_56 9.241569
Rin62_57 in62 in62_57 9.241569
Rin62_58 in62_57 in62_58 9.241569
Rin62_59 in62_58 in62_59 9.241569
Rin62_60 in62_59 in62_60 9.241569
Rin62_61 in62_60 in62_61 9.241569
Rin62_62 in62_61 in62_62 9.241569
Rin62_63 in62_62 in62_63 9.241569
Rin62_64 in62_63 in62_64 9.241569
Rin62_65 in62_64 in62_65 9.241569
Rin62_66 in62_65 in62_66 9.241569
Rin62_67 in62_66 in62_67 9.241569
Rin62_68 in62_67 in62_68 9.241569
Rin62_69 in62_68 in62_69 9.241569
Rin62_70 in62_69 in62_70 9.241569
Rin62_71 in62_70 in62_71 9.241569
Rin62_72 in62_71 in62_72 9.241569
Rin62_73 in62_72 in62_73 9.241569
Rin62_74 in62_73 in62_74 9.241569
Rin62_75 in62_74 in62_75 9.241569
Rin62_76 in62_75 in62_76 9.241569
Rin62_77 in62_76 in62_77 9.241569
Rin62_78 in62_77 in62_78 9.241569
Rin62_79 in62_78 in62_79 9.241569
Rin62_80 in62_79 in62_80 9.241569
Rin62_81 in62_80 in62_81 9.241569
Rin62_82 in62_81 in62_82 9.241569
Rin62_83 in62_82 in62_83 9.241569
Rin62_84 in62_83 in62_84 9.241569
Rin63_1 in63 in63_1 9.241569
Rin63_2 in63_1 in63_2 9.241569
Rin63_3 in63_2 in63_3 9.241569
Rin63_4 in63_3 in63_4 9.241569
Rin63_5 in63_4 in63_5 9.241569
Rin63_6 in63_5 in63_6 9.241569
Rin63_7 in63_6 in63_7 9.241569
Rin63_8 in63_7 in63_8 9.241569
Rin63_9 in63_8 in63_9 9.241569
Rin63_10 in63_9 in63_10 9.241569
Rin63_11 in63_10 in63_11 9.241569
Rin63_12 in63_11 in63_12 9.241569
Rin63_13 in63_12 in63_13 9.241569
Rin63_14 in63_13 in63_14 9.241569
Rin63_15 in63_14 in63_15 9.241569
Rin63_16 in63_15 in63_16 9.241569
Rin63_17 in63_16 in63_17 9.241569
Rin63_18 in63_17 in63_18 9.241569
Rin63_19 in63_18 in63_19 9.241569
Rin63_20 in63_19 in63_20 9.241569
Rin63_21 in63_20 in63_21 9.241569
Rin63_22 in63_21 in63_22 9.241569
Rin63_23 in63_22 in63_23 9.241569
Rin63_24 in63_23 in63_24 9.241569
Rin63_25 in63_24 in63_25 9.241569
Rin63_26 in63_25 in63_26 9.241569
Rin63_27 in63_26 in63_27 9.241569
Rin63_28 in63_27 in63_28 9.241569
Rin63_29 in63 in63_29 9.241569
Rin63_30 in63_29 in63_30 9.241569
Rin63_31 in63_30 in63_31 9.241569
Rin63_32 in63_31 in63_32 9.241569
Rin63_33 in63_32 in63_33 9.241569
Rin63_34 in63_33 in63_34 9.241569
Rin63_35 in63_34 in63_35 9.241569
Rin63_36 in63_35 in63_36 9.241569
Rin63_37 in63_36 in63_37 9.241569
Rin63_38 in63_37 in63_38 9.241569
Rin63_39 in63_38 in63_39 9.241569
Rin63_40 in63_39 in63_40 9.241569
Rin63_41 in63_40 in63_41 9.241569
Rin63_42 in63_41 in63_42 9.241569
Rin63_43 in63_42 in63_43 9.241569
Rin63_44 in63_43 in63_44 9.241569
Rin63_45 in63_44 in63_45 9.241569
Rin63_46 in63_45 in63_46 9.241569
Rin63_47 in63_46 in63_47 9.241569
Rin63_48 in63_47 in63_48 9.241569
Rin63_49 in63_48 in63_49 9.241569
Rin63_50 in63_49 in63_50 9.241569
Rin63_51 in63_50 in63_51 9.241569
Rin63_52 in63_51 in63_52 9.241569
Rin63_53 in63_52 in63_53 9.241569
Rin63_54 in63_53 in63_54 9.241569
Rin63_55 in63_54 in63_55 9.241569
Rin63_56 in63_55 in63_56 9.241569
Rin63_57 in63 in63_57 9.241569
Rin63_58 in63_57 in63_58 9.241569
Rin63_59 in63_58 in63_59 9.241569
Rin63_60 in63_59 in63_60 9.241569
Rin63_61 in63_60 in63_61 9.241569
Rin63_62 in63_61 in63_62 9.241569
Rin63_63 in63_62 in63_63 9.241569
Rin63_64 in63_63 in63_64 9.241569
Rin63_65 in63_64 in63_65 9.241569
Rin63_66 in63_65 in63_66 9.241569
Rin63_67 in63_66 in63_67 9.241569
Rin63_68 in63_67 in63_68 9.241569
Rin63_69 in63_68 in63_69 9.241569
Rin63_70 in63_69 in63_70 9.241569
Rin63_71 in63_70 in63_71 9.241569
Rin63_72 in63_71 in63_72 9.241569
Rin63_73 in63_72 in63_73 9.241569
Rin63_74 in63_73 in63_74 9.241569
Rin63_75 in63_74 in63_75 9.241569
Rin63_76 in63_75 in63_76 9.241569
Rin63_77 in63_76 in63_77 9.241569
Rin63_78 in63_77 in63_78 9.241569
Rin63_79 in63_78 in63_79 9.241569
Rin63_80 in63_79 in63_80 9.241569
Rin63_81 in63_80 in63_81 9.241569
Rin63_82 in63_81 in63_82 9.241569
Rin63_83 in63_82 in63_83 9.241569
Rin63_84 in63_83 in63_84 9.241569
Rin64_1 in64 in64_1 9.241569
Rin64_2 in64_1 in64_2 9.241569
Rin64_3 in64_2 in64_3 9.241569
Rin64_4 in64_3 in64_4 9.241569
Rin64_5 in64_4 in64_5 9.241569
Rin64_6 in64_5 in64_6 9.241569
Rin64_7 in64_6 in64_7 9.241569
Rin64_8 in64_7 in64_8 9.241569
Rin64_9 in64_8 in64_9 9.241569
Rin64_10 in64_9 in64_10 9.241569
Rin64_11 in64_10 in64_11 9.241569
Rin64_12 in64_11 in64_12 9.241569
Rin64_13 in64_12 in64_13 9.241569
Rin64_14 in64_13 in64_14 9.241569
Rin64_15 in64_14 in64_15 9.241569
Rin64_16 in64_15 in64_16 9.241569
Rin64_17 in64_16 in64_17 9.241569
Rin64_18 in64_17 in64_18 9.241569
Rin64_19 in64_18 in64_19 9.241569
Rin64_20 in64_19 in64_20 9.241569
Rin64_21 in64_20 in64_21 9.241569
Rin64_22 in64_21 in64_22 9.241569
Rin64_23 in64_22 in64_23 9.241569
Rin64_24 in64_23 in64_24 9.241569
Rin64_25 in64_24 in64_25 9.241569
Rin64_26 in64_25 in64_26 9.241569
Rin64_27 in64_26 in64_27 9.241569
Rin64_28 in64_27 in64_28 9.241569
Rin64_29 in64 in64_29 9.241569
Rin64_30 in64_29 in64_30 9.241569
Rin64_31 in64_30 in64_31 9.241569
Rin64_32 in64_31 in64_32 9.241569
Rin64_33 in64_32 in64_33 9.241569
Rin64_34 in64_33 in64_34 9.241569
Rin64_35 in64_34 in64_35 9.241569
Rin64_36 in64_35 in64_36 9.241569
Rin64_37 in64_36 in64_37 9.241569
Rin64_38 in64_37 in64_38 9.241569
Rin64_39 in64_38 in64_39 9.241569
Rin64_40 in64_39 in64_40 9.241569
Rin64_41 in64_40 in64_41 9.241569
Rin64_42 in64_41 in64_42 9.241569
Rin64_43 in64_42 in64_43 9.241569
Rin64_44 in64_43 in64_44 9.241569
Rin64_45 in64_44 in64_45 9.241569
Rin64_46 in64_45 in64_46 9.241569
Rin64_47 in64_46 in64_47 9.241569
Rin64_48 in64_47 in64_48 9.241569
Rin64_49 in64_48 in64_49 9.241569
Rin64_50 in64_49 in64_50 9.241569
Rin64_51 in64_50 in64_51 9.241569
Rin64_52 in64_51 in64_52 9.241569
Rin64_53 in64_52 in64_53 9.241569
Rin64_54 in64_53 in64_54 9.241569
Rin64_55 in64_54 in64_55 9.241569
Rin64_56 in64_55 in64_56 9.241569
Rin64_57 in64 in64_57 9.241569
Rin64_58 in64_57 in64_58 9.241569
Rin64_59 in64_58 in64_59 9.241569
Rin64_60 in64_59 in64_60 9.241569
Rin64_61 in64_60 in64_61 9.241569
Rin64_62 in64_61 in64_62 9.241569
Rin64_63 in64_62 in64_63 9.241569
Rin64_64 in64_63 in64_64 9.241569
Rin64_65 in64_64 in64_65 9.241569
Rin64_66 in64_65 in64_66 9.241569
Rin64_67 in64_66 in64_67 9.241569
Rin64_68 in64_67 in64_68 9.241569
Rin64_69 in64_68 in64_69 9.241569
Rin64_70 in64_69 in64_70 9.241569
Rin64_71 in64_70 in64_71 9.241569
Rin64_72 in64_71 in64_72 9.241569
Rin64_73 in64_72 in64_73 9.241569
Rin64_74 in64_73 in64_74 9.241569
Rin64_75 in64_74 in64_75 9.241569
Rin64_76 in64_75 in64_76 9.241569
Rin64_77 in64_76 in64_77 9.241569
Rin64_78 in64_77 in64_78 9.241569
Rin64_79 in64_78 in64_79 9.241569
Rin64_80 in64_79 in64_80 9.241569
Rin64_81 in64_80 in64_81 9.241569
Rin64_82 in64_81 in64_82 9.241569
Rin64_83 in64_82 in64_83 9.241569
Rin64_84 in64_83 in64_84 9.241569
Rin65_1 in65 in65_1 9.241569
Rin65_2 in65_1 in65_2 9.241569
Rin65_3 in65_2 in65_3 9.241569
Rin65_4 in65_3 in65_4 9.241569
Rin65_5 in65_4 in65_5 9.241569
Rin65_6 in65_5 in65_6 9.241569
Rin65_7 in65_6 in65_7 9.241569
Rin65_8 in65_7 in65_8 9.241569
Rin65_9 in65_8 in65_9 9.241569
Rin65_10 in65_9 in65_10 9.241569
Rin65_11 in65_10 in65_11 9.241569
Rin65_12 in65_11 in65_12 9.241569
Rin65_13 in65_12 in65_13 9.241569
Rin65_14 in65_13 in65_14 9.241569
Rin65_15 in65_14 in65_15 9.241569
Rin65_16 in65_15 in65_16 9.241569
Rin65_17 in65_16 in65_17 9.241569
Rin65_18 in65_17 in65_18 9.241569
Rin65_19 in65_18 in65_19 9.241569
Rin65_20 in65_19 in65_20 9.241569
Rin65_21 in65_20 in65_21 9.241569
Rin65_22 in65_21 in65_22 9.241569
Rin65_23 in65_22 in65_23 9.241569
Rin65_24 in65_23 in65_24 9.241569
Rin65_25 in65_24 in65_25 9.241569
Rin65_26 in65_25 in65_26 9.241569
Rin65_27 in65_26 in65_27 9.241569
Rin65_28 in65_27 in65_28 9.241569
Rin65_29 in65 in65_29 9.241569
Rin65_30 in65_29 in65_30 9.241569
Rin65_31 in65_30 in65_31 9.241569
Rin65_32 in65_31 in65_32 9.241569
Rin65_33 in65_32 in65_33 9.241569
Rin65_34 in65_33 in65_34 9.241569
Rin65_35 in65_34 in65_35 9.241569
Rin65_36 in65_35 in65_36 9.241569
Rin65_37 in65_36 in65_37 9.241569
Rin65_38 in65_37 in65_38 9.241569
Rin65_39 in65_38 in65_39 9.241569
Rin65_40 in65_39 in65_40 9.241569
Rin65_41 in65_40 in65_41 9.241569
Rin65_42 in65_41 in65_42 9.241569
Rin65_43 in65_42 in65_43 9.241569
Rin65_44 in65_43 in65_44 9.241569
Rin65_45 in65_44 in65_45 9.241569
Rin65_46 in65_45 in65_46 9.241569
Rin65_47 in65_46 in65_47 9.241569
Rin65_48 in65_47 in65_48 9.241569
Rin65_49 in65_48 in65_49 9.241569
Rin65_50 in65_49 in65_50 9.241569
Rin65_51 in65_50 in65_51 9.241569
Rin65_52 in65_51 in65_52 9.241569
Rin65_53 in65_52 in65_53 9.241569
Rin65_54 in65_53 in65_54 9.241569
Rin65_55 in65_54 in65_55 9.241569
Rin65_56 in65_55 in65_56 9.241569
Rin65_57 in65 in65_57 9.241569
Rin65_58 in65_57 in65_58 9.241569
Rin65_59 in65_58 in65_59 9.241569
Rin65_60 in65_59 in65_60 9.241569
Rin65_61 in65_60 in65_61 9.241569
Rin65_62 in65_61 in65_62 9.241569
Rin65_63 in65_62 in65_63 9.241569
Rin65_64 in65_63 in65_64 9.241569
Rin65_65 in65_64 in65_65 9.241569
Rin65_66 in65_65 in65_66 9.241569
Rin65_67 in65_66 in65_67 9.241569
Rin65_68 in65_67 in65_68 9.241569
Rin65_69 in65_68 in65_69 9.241569
Rin65_70 in65_69 in65_70 9.241569
Rin65_71 in65_70 in65_71 9.241569
Rin65_72 in65_71 in65_72 9.241569
Rin65_73 in65_72 in65_73 9.241569
Rin65_74 in65_73 in65_74 9.241569
Rin65_75 in65_74 in65_75 9.241569
Rin65_76 in65_75 in65_76 9.241569
Rin65_77 in65_76 in65_77 9.241569
Rin65_78 in65_77 in65_78 9.241569
Rin65_79 in65_78 in65_79 9.241569
Rin65_80 in65_79 in65_80 9.241569
Rin65_81 in65_80 in65_81 9.241569
Rin65_82 in65_81 in65_82 9.241569
Rin65_83 in65_82 in65_83 9.241569
Rin65_84 in65_83 in65_84 9.241569
Rin66_1 in66 in66_1 9.241569
Rin66_2 in66_1 in66_2 9.241569
Rin66_3 in66_2 in66_3 9.241569
Rin66_4 in66_3 in66_4 9.241569
Rin66_5 in66_4 in66_5 9.241569
Rin66_6 in66_5 in66_6 9.241569
Rin66_7 in66_6 in66_7 9.241569
Rin66_8 in66_7 in66_8 9.241569
Rin66_9 in66_8 in66_9 9.241569
Rin66_10 in66_9 in66_10 9.241569
Rin66_11 in66_10 in66_11 9.241569
Rin66_12 in66_11 in66_12 9.241569
Rin66_13 in66_12 in66_13 9.241569
Rin66_14 in66_13 in66_14 9.241569
Rin66_15 in66_14 in66_15 9.241569
Rin66_16 in66_15 in66_16 9.241569
Rin66_17 in66_16 in66_17 9.241569
Rin66_18 in66_17 in66_18 9.241569
Rin66_19 in66_18 in66_19 9.241569
Rin66_20 in66_19 in66_20 9.241569
Rin66_21 in66_20 in66_21 9.241569
Rin66_22 in66_21 in66_22 9.241569
Rin66_23 in66_22 in66_23 9.241569
Rin66_24 in66_23 in66_24 9.241569
Rin66_25 in66_24 in66_25 9.241569
Rin66_26 in66_25 in66_26 9.241569
Rin66_27 in66_26 in66_27 9.241569
Rin66_28 in66_27 in66_28 9.241569
Rin66_29 in66 in66_29 9.241569
Rin66_30 in66_29 in66_30 9.241569
Rin66_31 in66_30 in66_31 9.241569
Rin66_32 in66_31 in66_32 9.241569
Rin66_33 in66_32 in66_33 9.241569
Rin66_34 in66_33 in66_34 9.241569
Rin66_35 in66_34 in66_35 9.241569
Rin66_36 in66_35 in66_36 9.241569
Rin66_37 in66_36 in66_37 9.241569
Rin66_38 in66_37 in66_38 9.241569
Rin66_39 in66_38 in66_39 9.241569
Rin66_40 in66_39 in66_40 9.241569
Rin66_41 in66_40 in66_41 9.241569
Rin66_42 in66_41 in66_42 9.241569
Rin66_43 in66_42 in66_43 9.241569
Rin66_44 in66_43 in66_44 9.241569
Rin66_45 in66_44 in66_45 9.241569
Rin66_46 in66_45 in66_46 9.241569
Rin66_47 in66_46 in66_47 9.241569
Rin66_48 in66_47 in66_48 9.241569
Rin66_49 in66_48 in66_49 9.241569
Rin66_50 in66_49 in66_50 9.241569
Rin66_51 in66_50 in66_51 9.241569
Rin66_52 in66_51 in66_52 9.241569
Rin66_53 in66_52 in66_53 9.241569
Rin66_54 in66_53 in66_54 9.241569
Rin66_55 in66_54 in66_55 9.241569
Rin66_56 in66_55 in66_56 9.241569
Rin66_57 in66 in66_57 9.241569
Rin66_58 in66_57 in66_58 9.241569
Rin66_59 in66_58 in66_59 9.241569
Rin66_60 in66_59 in66_60 9.241569
Rin66_61 in66_60 in66_61 9.241569
Rin66_62 in66_61 in66_62 9.241569
Rin66_63 in66_62 in66_63 9.241569
Rin66_64 in66_63 in66_64 9.241569
Rin66_65 in66_64 in66_65 9.241569
Rin66_66 in66_65 in66_66 9.241569
Rin66_67 in66_66 in66_67 9.241569
Rin66_68 in66_67 in66_68 9.241569
Rin66_69 in66_68 in66_69 9.241569
Rin66_70 in66_69 in66_70 9.241569
Rin66_71 in66_70 in66_71 9.241569
Rin66_72 in66_71 in66_72 9.241569
Rin66_73 in66_72 in66_73 9.241569
Rin66_74 in66_73 in66_74 9.241569
Rin66_75 in66_74 in66_75 9.241569
Rin66_76 in66_75 in66_76 9.241569
Rin66_77 in66_76 in66_77 9.241569
Rin66_78 in66_77 in66_78 9.241569
Rin66_79 in66_78 in66_79 9.241569
Rin66_80 in66_79 in66_80 9.241569
Rin66_81 in66_80 in66_81 9.241569
Rin66_82 in66_81 in66_82 9.241569
Rin66_83 in66_82 in66_83 9.241569
Rin66_84 in66_83 in66_84 9.241569
Rin67_1 in67 in67_1 9.241569
Rin67_2 in67_1 in67_2 9.241569
Rin67_3 in67_2 in67_3 9.241569
Rin67_4 in67_3 in67_4 9.241569
Rin67_5 in67_4 in67_5 9.241569
Rin67_6 in67_5 in67_6 9.241569
Rin67_7 in67_6 in67_7 9.241569
Rin67_8 in67_7 in67_8 9.241569
Rin67_9 in67_8 in67_9 9.241569
Rin67_10 in67_9 in67_10 9.241569
Rin67_11 in67_10 in67_11 9.241569
Rin67_12 in67_11 in67_12 9.241569
Rin67_13 in67_12 in67_13 9.241569
Rin67_14 in67_13 in67_14 9.241569
Rin67_15 in67_14 in67_15 9.241569
Rin67_16 in67_15 in67_16 9.241569
Rin67_17 in67_16 in67_17 9.241569
Rin67_18 in67_17 in67_18 9.241569
Rin67_19 in67_18 in67_19 9.241569
Rin67_20 in67_19 in67_20 9.241569
Rin67_21 in67_20 in67_21 9.241569
Rin67_22 in67_21 in67_22 9.241569
Rin67_23 in67_22 in67_23 9.241569
Rin67_24 in67_23 in67_24 9.241569
Rin67_25 in67_24 in67_25 9.241569
Rin67_26 in67_25 in67_26 9.241569
Rin67_27 in67_26 in67_27 9.241569
Rin67_28 in67_27 in67_28 9.241569
Rin67_29 in67 in67_29 9.241569
Rin67_30 in67_29 in67_30 9.241569
Rin67_31 in67_30 in67_31 9.241569
Rin67_32 in67_31 in67_32 9.241569
Rin67_33 in67_32 in67_33 9.241569
Rin67_34 in67_33 in67_34 9.241569
Rin67_35 in67_34 in67_35 9.241569
Rin67_36 in67_35 in67_36 9.241569
Rin67_37 in67_36 in67_37 9.241569
Rin67_38 in67_37 in67_38 9.241569
Rin67_39 in67_38 in67_39 9.241569
Rin67_40 in67_39 in67_40 9.241569
Rin67_41 in67_40 in67_41 9.241569
Rin67_42 in67_41 in67_42 9.241569
Rin67_43 in67_42 in67_43 9.241569
Rin67_44 in67_43 in67_44 9.241569
Rin67_45 in67_44 in67_45 9.241569
Rin67_46 in67_45 in67_46 9.241569
Rin67_47 in67_46 in67_47 9.241569
Rin67_48 in67_47 in67_48 9.241569
Rin67_49 in67_48 in67_49 9.241569
Rin67_50 in67_49 in67_50 9.241569
Rin67_51 in67_50 in67_51 9.241569
Rin67_52 in67_51 in67_52 9.241569
Rin67_53 in67_52 in67_53 9.241569
Rin67_54 in67_53 in67_54 9.241569
Rin67_55 in67_54 in67_55 9.241569
Rin67_56 in67_55 in67_56 9.241569
Rin67_57 in67 in67_57 9.241569
Rin67_58 in67_57 in67_58 9.241569
Rin67_59 in67_58 in67_59 9.241569
Rin67_60 in67_59 in67_60 9.241569
Rin67_61 in67_60 in67_61 9.241569
Rin67_62 in67_61 in67_62 9.241569
Rin67_63 in67_62 in67_63 9.241569
Rin67_64 in67_63 in67_64 9.241569
Rin67_65 in67_64 in67_65 9.241569
Rin67_66 in67_65 in67_66 9.241569
Rin67_67 in67_66 in67_67 9.241569
Rin67_68 in67_67 in67_68 9.241569
Rin67_69 in67_68 in67_69 9.241569
Rin67_70 in67_69 in67_70 9.241569
Rin67_71 in67_70 in67_71 9.241569
Rin67_72 in67_71 in67_72 9.241569
Rin67_73 in67_72 in67_73 9.241569
Rin67_74 in67_73 in67_74 9.241569
Rin67_75 in67_74 in67_75 9.241569
Rin67_76 in67_75 in67_76 9.241569
Rin67_77 in67_76 in67_77 9.241569
Rin67_78 in67_77 in67_78 9.241569
Rin67_79 in67_78 in67_79 9.241569
Rin67_80 in67_79 in67_80 9.241569
Rin67_81 in67_80 in67_81 9.241569
Rin67_82 in67_81 in67_82 9.241569
Rin67_83 in67_82 in67_83 9.241569
Rin67_84 in67_83 in67_84 9.241569
Rin68_1 in68 in68_1 9.241569
Rin68_2 in68_1 in68_2 9.241569
Rin68_3 in68_2 in68_3 9.241569
Rin68_4 in68_3 in68_4 9.241569
Rin68_5 in68_4 in68_5 9.241569
Rin68_6 in68_5 in68_6 9.241569
Rin68_7 in68_6 in68_7 9.241569
Rin68_8 in68_7 in68_8 9.241569
Rin68_9 in68_8 in68_9 9.241569
Rin68_10 in68_9 in68_10 9.241569
Rin68_11 in68_10 in68_11 9.241569
Rin68_12 in68_11 in68_12 9.241569
Rin68_13 in68_12 in68_13 9.241569
Rin68_14 in68_13 in68_14 9.241569
Rin68_15 in68_14 in68_15 9.241569
Rin68_16 in68_15 in68_16 9.241569
Rin68_17 in68_16 in68_17 9.241569
Rin68_18 in68_17 in68_18 9.241569
Rin68_19 in68_18 in68_19 9.241569
Rin68_20 in68_19 in68_20 9.241569
Rin68_21 in68_20 in68_21 9.241569
Rin68_22 in68_21 in68_22 9.241569
Rin68_23 in68_22 in68_23 9.241569
Rin68_24 in68_23 in68_24 9.241569
Rin68_25 in68_24 in68_25 9.241569
Rin68_26 in68_25 in68_26 9.241569
Rin68_27 in68_26 in68_27 9.241569
Rin68_28 in68_27 in68_28 9.241569
Rin68_29 in68 in68_29 9.241569
Rin68_30 in68_29 in68_30 9.241569
Rin68_31 in68_30 in68_31 9.241569
Rin68_32 in68_31 in68_32 9.241569
Rin68_33 in68_32 in68_33 9.241569
Rin68_34 in68_33 in68_34 9.241569
Rin68_35 in68_34 in68_35 9.241569
Rin68_36 in68_35 in68_36 9.241569
Rin68_37 in68_36 in68_37 9.241569
Rin68_38 in68_37 in68_38 9.241569
Rin68_39 in68_38 in68_39 9.241569
Rin68_40 in68_39 in68_40 9.241569
Rin68_41 in68_40 in68_41 9.241569
Rin68_42 in68_41 in68_42 9.241569
Rin68_43 in68_42 in68_43 9.241569
Rin68_44 in68_43 in68_44 9.241569
Rin68_45 in68_44 in68_45 9.241569
Rin68_46 in68_45 in68_46 9.241569
Rin68_47 in68_46 in68_47 9.241569
Rin68_48 in68_47 in68_48 9.241569
Rin68_49 in68_48 in68_49 9.241569
Rin68_50 in68_49 in68_50 9.241569
Rin68_51 in68_50 in68_51 9.241569
Rin68_52 in68_51 in68_52 9.241569
Rin68_53 in68_52 in68_53 9.241569
Rin68_54 in68_53 in68_54 9.241569
Rin68_55 in68_54 in68_55 9.241569
Rin68_56 in68_55 in68_56 9.241569
Rin68_57 in68 in68_57 9.241569
Rin68_58 in68_57 in68_58 9.241569
Rin68_59 in68_58 in68_59 9.241569
Rin68_60 in68_59 in68_60 9.241569
Rin68_61 in68_60 in68_61 9.241569
Rin68_62 in68_61 in68_62 9.241569
Rin68_63 in68_62 in68_63 9.241569
Rin68_64 in68_63 in68_64 9.241569
Rin68_65 in68_64 in68_65 9.241569
Rin68_66 in68_65 in68_66 9.241569
Rin68_67 in68_66 in68_67 9.241569
Rin68_68 in68_67 in68_68 9.241569
Rin68_69 in68_68 in68_69 9.241569
Rin68_70 in68_69 in68_70 9.241569
Rin68_71 in68_70 in68_71 9.241569
Rin68_72 in68_71 in68_72 9.241569
Rin68_73 in68_72 in68_73 9.241569
Rin68_74 in68_73 in68_74 9.241569
Rin68_75 in68_74 in68_75 9.241569
Rin68_76 in68_75 in68_76 9.241569
Rin68_77 in68_76 in68_77 9.241569
Rin68_78 in68_77 in68_78 9.241569
Rin68_79 in68_78 in68_79 9.241569
Rin68_80 in68_79 in68_80 9.241569
Rin68_81 in68_80 in68_81 9.241569
Rin68_82 in68_81 in68_82 9.241569
Rin68_83 in68_82 in68_83 9.241569
Rin68_84 in68_83 in68_84 9.241569
Rin69_1 in69 in69_1 9.241569
Rin69_2 in69_1 in69_2 9.241569
Rin69_3 in69_2 in69_3 9.241569
Rin69_4 in69_3 in69_4 9.241569
Rin69_5 in69_4 in69_5 9.241569
Rin69_6 in69_5 in69_6 9.241569
Rin69_7 in69_6 in69_7 9.241569
Rin69_8 in69_7 in69_8 9.241569
Rin69_9 in69_8 in69_9 9.241569
Rin69_10 in69_9 in69_10 9.241569
Rin69_11 in69_10 in69_11 9.241569
Rin69_12 in69_11 in69_12 9.241569
Rin69_13 in69_12 in69_13 9.241569
Rin69_14 in69_13 in69_14 9.241569
Rin69_15 in69_14 in69_15 9.241569
Rin69_16 in69_15 in69_16 9.241569
Rin69_17 in69_16 in69_17 9.241569
Rin69_18 in69_17 in69_18 9.241569
Rin69_19 in69_18 in69_19 9.241569
Rin69_20 in69_19 in69_20 9.241569
Rin69_21 in69_20 in69_21 9.241569
Rin69_22 in69_21 in69_22 9.241569
Rin69_23 in69_22 in69_23 9.241569
Rin69_24 in69_23 in69_24 9.241569
Rin69_25 in69_24 in69_25 9.241569
Rin69_26 in69_25 in69_26 9.241569
Rin69_27 in69_26 in69_27 9.241569
Rin69_28 in69_27 in69_28 9.241569
Rin69_29 in69 in69_29 9.241569
Rin69_30 in69_29 in69_30 9.241569
Rin69_31 in69_30 in69_31 9.241569
Rin69_32 in69_31 in69_32 9.241569
Rin69_33 in69_32 in69_33 9.241569
Rin69_34 in69_33 in69_34 9.241569
Rin69_35 in69_34 in69_35 9.241569
Rin69_36 in69_35 in69_36 9.241569
Rin69_37 in69_36 in69_37 9.241569
Rin69_38 in69_37 in69_38 9.241569
Rin69_39 in69_38 in69_39 9.241569
Rin69_40 in69_39 in69_40 9.241569
Rin69_41 in69_40 in69_41 9.241569
Rin69_42 in69_41 in69_42 9.241569
Rin69_43 in69_42 in69_43 9.241569
Rin69_44 in69_43 in69_44 9.241569
Rin69_45 in69_44 in69_45 9.241569
Rin69_46 in69_45 in69_46 9.241569
Rin69_47 in69_46 in69_47 9.241569
Rin69_48 in69_47 in69_48 9.241569
Rin69_49 in69_48 in69_49 9.241569
Rin69_50 in69_49 in69_50 9.241569
Rin69_51 in69_50 in69_51 9.241569
Rin69_52 in69_51 in69_52 9.241569
Rin69_53 in69_52 in69_53 9.241569
Rin69_54 in69_53 in69_54 9.241569
Rin69_55 in69_54 in69_55 9.241569
Rin69_56 in69_55 in69_56 9.241569
Rin69_57 in69 in69_57 9.241569
Rin69_58 in69_57 in69_58 9.241569
Rin69_59 in69_58 in69_59 9.241569
Rin69_60 in69_59 in69_60 9.241569
Rin69_61 in69_60 in69_61 9.241569
Rin69_62 in69_61 in69_62 9.241569
Rin69_63 in69_62 in69_63 9.241569
Rin69_64 in69_63 in69_64 9.241569
Rin69_65 in69_64 in69_65 9.241569
Rin69_66 in69_65 in69_66 9.241569
Rin69_67 in69_66 in69_67 9.241569
Rin69_68 in69_67 in69_68 9.241569
Rin69_69 in69_68 in69_69 9.241569
Rin69_70 in69_69 in69_70 9.241569
Rin69_71 in69_70 in69_71 9.241569
Rin69_72 in69_71 in69_72 9.241569
Rin69_73 in69_72 in69_73 9.241569
Rin69_74 in69_73 in69_74 9.241569
Rin69_75 in69_74 in69_75 9.241569
Rin69_76 in69_75 in69_76 9.241569
Rin69_77 in69_76 in69_77 9.241569
Rin69_78 in69_77 in69_78 9.241569
Rin69_79 in69_78 in69_79 9.241569
Rin69_80 in69_79 in69_80 9.241569
Rin69_81 in69_80 in69_81 9.241569
Rin69_82 in69_81 in69_82 9.241569
Rin69_83 in69_82 in69_83 9.241569
Rin69_84 in69_83 in69_84 9.241569
Rin70_1 in70 in70_1 9.241569
Rin70_2 in70_1 in70_2 9.241569
Rin70_3 in70_2 in70_3 9.241569
Rin70_4 in70_3 in70_4 9.241569
Rin70_5 in70_4 in70_5 9.241569
Rin70_6 in70_5 in70_6 9.241569
Rin70_7 in70_6 in70_7 9.241569
Rin70_8 in70_7 in70_8 9.241569
Rin70_9 in70_8 in70_9 9.241569
Rin70_10 in70_9 in70_10 9.241569
Rin70_11 in70_10 in70_11 9.241569
Rin70_12 in70_11 in70_12 9.241569
Rin70_13 in70_12 in70_13 9.241569
Rin70_14 in70_13 in70_14 9.241569
Rin70_15 in70_14 in70_15 9.241569
Rin70_16 in70_15 in70_16 9.241569
Rin70_17 in70_16 in70_17 9.241569
Rin70_18 in70_17 in70_18 9.241569
Rin70_19 in70_18 in70_19 9.241569
Rin70_20 in70_19 in70_20 9.241569
Rin70_21 in70_20 in70_21 9.241569
Rin70_22 in70_21 in70_22 9.241569
Rin70_23 in70_22 in70_23 9.241569
Rin70_24 in70_23 in70_24 9.241569
Rin70_25 in70_24 in70_25 9.241569
Rin70_26 in70_25 in70_26 9.241569
Rin70_27 in70_26 in70_27 9.241569
Rin70_28 in70_27 in70_28 9.241569
Rin70_29 in70 in70_29 9.241569
Rin70_30 in70_29 in70_30 9.241569
Rin70_31 in70_30 in70_31 9.241569
Rin70_32 in70_31 in70_32 9.241569
Rin70_33 in70_32 in70_33 9.241569
Rin70_34 in70_33 in70_34 9.241569
Rin70_35 in70_34 in70_35 9.241569
Rin70_36 in70_35 in70_36 9.241569
Rin70_37 in70_36 in70_37 9.241569
Rin70_38 in70_37 in70_38 9.241569
Rin70_39 in70_38 in70_39 9.241569
Rin70_40 in70_39 in70_40 9.241569
Rin70_41 in70_40 in70_41 9.241569
Rin70_42 in70_41 in70_42 9.241569
Rin70_43 in70_42 in70_43 9.241569
Rin70_44 in70_43 in70_44 9.241569
Rin70_45 in70_44 in70_45 9.241569
Rin70_46 in70_45 in70_46 9.241569
Rin70_47 in70_46 in70_47 9.241569
Rin70_48 in70_47 in70_48 9.241569
Rin70_49 in70_48 in70_49 9.241569
Rin70_50 in70_49 in70_50 9.241569
Rin70_51 in70_50 in70_51 9.241569
Rin70_52 in70_51 in70_52 9.241569
Rin70_53 in70_52 in70_53 9.241569
Rin70_54 in70_53 in70_54 9.241569
Rin70_55 in70_54 in70_55 9.241569
Rin70_56 in70_55 in70_56 9.241569
Rin70_57 in70 in70_57 9.241569
Rin70_58 in70_57 in70_58 9.241569
Rin70_59 in70_58 in70_59 9.241569
Rin70_60 in70_59 in70_60 9.241569
Rin70_61 in70_60 in70_61 9.241569
Rin70_62 in70_61 in70_62 9.241569
Rin70_63 in70_62 in70_63 9.241569
Rin70_64 in70_63 in70_64 9.241569
Rin70_65 in70_64 in70_65 9.241569
Rin70_66 in70_65 in70_66 9.241569
Rin70_67 in70_66 in70_67 9.241569
Rin70_68 in70_67 in70_68 9.241569
Rin70_69 in70_68 in70_69 9.241569
Rin70_70 in70_69 in70_70 9.241569
Rin70_71 in70_70 in70_71 9.241569
Rin70_72 in70_71 in70_72 9.241569
Rin70_73 in70_72 in70_73 9.241569
Rin70_74 in70_73 in70_74 9.241569
Rin70_75 in70_74 in70_75 9.241569
Rin70_76 in70_75 in70_76 9.241569
Rin70_77 in70_76 in70_77 9.241569
Rin70_78 in70_77 in70_78 9.241569
Rin70_79 in70_78 in70_79 9.241569
Rin70_80 in70_79 in70_80 9.241569
Rin70_81 in70_80 in70_81 9.241569
Rin70_82 in70_81 in70_82 9.241569
Rin70_83 in70_82 in70_83 9.241569
Rin70_84 in70_83 in70_84 9.241569
Rin71_1 in71 in71_1 9.241569
Rin71_2 in71_1 in71_2 9.241569
Rin71_3 in71_2 in71_3 9.241569
Rin71_4 in71_3 in71_4 9.241569
Rin71_5 in71_4 in71_5 9.241569
Rin71_6 in71_5 in71_6 9.241569
Rin71_7 in71_6 in71_7 9.241569
Rin71_8 in71_7 in71_8 9.241569
Rin71_9 in71_8 in71_9 9.241569
Rin71_10 in71_9 in71_10 9.241569
Rin71_11 in71_10 in71_11 9.241569
Rin71_12 in71_11 in71_12 9.241569
Rin71_13 in71_12 in71_13 9.241569
Rin71_14 in71_13 in71_14 9.241569
Rin71_15 in71_14 in71_15 9.241569
Rin71_16 in71_15 in71_16 9.241569
Rin71_17 in71_16 in71_17 9.241569
Rin71_18 in71_17 in71_18 9.241569
Rin71_19 in71_18 in71_19 9.241569
Rin71_20 in71_19 in71_20 9.241569
Rin71_21 in71_20 in71_21 9.241569
Rin71_22 in71_21 in71_22 9.241569
Rin71_23 in71_22 in71_23 9.241569
Rin71_24 in71_23 in71_24 9.241569
Rin71_25 in71_24 in71_25 9.241569
Rin71_26 in71_25 in71_26 9.241569
Rin71_27 in71_26 in71_27 9.241569
Rin71_28 in71_27 in71_28 9.241569
Rin71_29 in71 in71_29 9.241569
Rin71_30 in71_29 in71_30 9.241569
Rin71_31 in71_30 in71_31 9.241569
Rin71_32 in71_31 in71_32 9.241569
Rin71_33 in71_32 in71_33 9.241569
Rin71_34 in71_33 in71_34 9.241569
Rin71_35 in71_34 in71_35 9.241569
Rin71_36 in71_35 in71_36 9.241569
Rin71_37 in71_36 in71_37 9.241569
Rin71_38 in71_37 in71_38 9.241569
Rin71_39 in71_38 in71_39 9.241569
Rin71_40 in71_39 in71_40 9.241569
Rin71_41 in71_40 in71_41 9.241569
Rin71_42 in71_41 in71_42 9.241569
Rin71_43 in71_42 in71_43 9.241569
Rin71_44 in71_43 in71_44 9.241569
Rin71_45 in71_44 in71_45 9.241569
Rin71_46 in71_45 in71_46 9.241569
Rin71_47 in71_46 in71_47 9.241569
Rin71_48 in71_47 in71_48 9.241569
Rin71_49 in71_48 in71_49 9.241569
Rin71_50 in71_49 in71_50 9.241569
Rin71_51 in71_50 in71_51 9.241569
Rin71_52 in71_51 in71_52 9.241569
Rin71_53 in71_52 in71_53 9.241569
Rin71_54 in71_53 in71_54 9.241569
Rin71_55 in71_54 in71_55 9.241569
Rin71_56 in71_55 in71_56 9.241569
Rin71_57 in71 in71_57 9.241569
Rin71_58 in71_57 in71_58 9.241569
Rin71_59 in71_58 in71_59 9.241569
Rin71_60 in71_59 in71_60 9.241569
Rin71_61 in71_60 in71_61 9.241569
Rin71_62 in71_61 in71_62 9.241569
Rin71_63 in71_62 in71_63 9.241569
Rin71_64 in71_63 in71_64 9.241569
Rin71_65 in71_64 in71_65 9.241569
Rin71_66 in71_65 in71_66 9.241569
Rin71_67 in71_66 in71_67 9.241569
Rin71_68 in71_67 in71_68 9.241569
Rin71_69 in71_68 in71_69 9.241569
Rin71_70 in71_69 in71_70 9.241569
Rin71_71 in71_70 in71_71 9.241569
Rin71_72 in71_71 in71_72 9.241569
Rin71_73 in71_72 in71_73 9.241569
Rin71_74 in71_73 in71_74 9.241569
Rin71_75 in71_74 in71_75 9.241569
Rin71_76 in71_75 in71_76 9.241569
Rin71_77 in71_76 in71_77 9.241569
Rin71_78 in71_77 in71_78 9.241569
Rin71_79 in71_78 in71_79 9.241569
Rin71_80 in71_79 in71_80 9.241569
Rin71_81 in71_80 in71_81 9.241569
Rin71_82 in71_81 in71_82 9.241569
Rin71_83 in71_82 in71_83 9.241569
Rin71_84 in71_83 in71_84 9.241569
Rin72_1 in72 in72_1 9.241569
Rin72_2 in72_1 in72_2 9.241569
Rin72_3 in72_2 in72_3 9.241569
Rin72_4 in72_3 in72_4 9.241569
Rin72_5 in72_4 in72_5 9.241569
Rin72_6 in72_5 in72_6 9.241569
Rin72_7 in72_6 in72_7 9.241569
Rin72_8 in72_7 in72_8 9.241569
Rin72_9 in72_8 in72_9 9.241569
Rin72_10 in72_9 in72_10 9.241569
Rin72_11 in72_10 in72_11 9.241569
Rin72_12 in72_11 in72_12 9.241569
Rin72_13 in72_12 in72_13 9.241569
Rin72_14 in72_13 in72_14 9.241569
Rin72_15 in72_14 in72_15 9.241569
Rin72_16 in72_15 in72_16 9.241569
Rin72_17 in72_16 in72_17 9.241569
Rin72_18 in72_17 in72_18 9.241569
Rin72_19 in72_18 in72_19 9.241569
Rin72_20 in72_19 in72_20 9.241569
Rin72_21 in72_20 in72_21 9.241569
Rin72_22 in72_21 in72_22 9.241569
Rin72_23 in72_22 in72_23 9.241569
Rin72_24 in72_23 in72_24 9.241569
Rin72_25 in72_24 in72_25 9.241569
Rin72_26 in72_25 in72_26 9.241569
Rin72_27 in72_26 in72_27 9.241569
Rin72_28 in72_27 in72_28 9.241569
Rin72_29 in72 in72_29 9.241569
Rin72_30 in72_29 in72_30 9.241569
Rin72_31 in72_30 in72_31 9.241569
Rin72_32 in72_31 in72_32 9.241569
Rin72_33 in72_32 in72_33 9.241569
Rin72_34 in72_33 in72_34 9.241569
Rin72_35 in72_34 in72_35 9.241569
Rin72_36 in72_35 in72_36 9.241569
Rin72_37 in72_36 in72_37 9.241569
Rin72_38 in72_37 in72_38 9.241569
Rin72_39 in72_38 in72_39 9.241569
Rin72_40 in72_39 in72_40 9.241569
Rin72_41 in72_40 in72_41 9.241569
Rin72_42 in72_41 in72_42 9.241569
Rin72_43 in72_42 in72_43 9.241569
Rin72_44 in72_43 in72_44 9.241569
Rin72_45 in72_44 in72_45 9.241569
Rin72_46 in72_45 in72_46 9.241569
Rin72_47 in72_46 in72_47 9.241569
Rin72_48 in72_47 in72_48 9.241569
Rin72_49 in72_48 in72_49 9.241569
Rin72_50 in72_49 in72_50 9.241569
Rin72_51 in72_50 in72_51 9.241569
Rin72_52 in72_51 in72_52 9.241569
Rin72_53 in72_52 in72_53 9.241569
Rin72_54 in72_53 in72_54 9.241569
Rin72_55 in72_54 in72_55 9.241569
Rin72_56 in72_55 in72_56 9.241569
Rin72_57 in72 in72_57 9.241569
Rin72_58 in72_57 in72_58 9.241569
Rin72_59 in72_58 in72_59 9.241569
Rin72_60 in72_59 in72_60 9.241569
Rin72_61 in72_60 in72_61 9.241569
Rin72_62 in72_61 in72_62 9.241569
Rin72_63 in72_62 in72_63 9.241569
Rin72_64 in72_63 in72_64 9.241569
Rin72_65 in72_64 in72_65 9.241569
Rin72_66 in72_65 in72_66 9.241569
Rin72_67 in72_66 in72_67 9.241569
Rin72_68 in72_67 in72_68 9.241569
Rin72_69 in72_68 in72_69 9.241569
Rin72_70 in72_69 in72_70 9.241569
Rin72_71 in72_70 in72_71 9.241569
Rin72_72 in72_71 in72_72 9.241569
Rin72_73 in72_72 in72_73 9.241569
Rin72_74 in72_73 in72_74 9.241569
Rin72_75 in72_74 in72_75 9.241569
Rin72_76 in72_75 in72_76 9.241569
Rin72_77 in72_76 in72_77 9.241569
Rin72_78 in72_77 in72_78 9.241569
Rin72_79 in72_78 in72_79 9.241569
Rin72_80 in72_79 in72_80 9.241569
Rin72_81 in72_80 in72_81 9.241569
Rin72_82 in72_81 in72_82 9.241569
Rin72_83 in72_82 in72_83 9.241569
Rin72_84 in72_83 in72_84 9.241569
Rin73_1 in73 in73_1 9.241569
Rin73_2 in73_1 in73_2 9.241569
Rin73_3 in73_2 in73_3 9.241569
Rin73_4 in73_3 in73_4 9.241569
Rin73_5 in73_4 in73_5 9.241569
Rin73_6 in73_5 in73_6 9.241569
Rin73_7 in73_6 in73_7 9.241569
Rin73_8 in73_7 in73_8 9.241569
Rin73_9 in73_8 in73_9 9.241569
Rin73_10 in73_9 in73_10 9.241569
Rin73_11 in73_10 in73_11 9.241569
Rin73_12 in73_11 in73_12 9.241569
Rin73_13 in73_12 in73_13 9.241569
Rin73_14 in73_13 in73_14 9.241569
Rin73_15 in73_14 in73_15 9.241569
Rin73_16 in73_15 in73_16 9.241569
Rin73_17 in73_16 in73_17 9.241569
Rin73_18 in73_17 in73_18 9.241569
Rin73_19 in73_18 in73_19 9.241569
Rin73_20 in73_19 in73_20 9.241569
Rin73_21 in73_20 in73_21 9.241569
Rin73_22 in73_21 in73_22 9.241569
Rin73_23 in73_22 in73_23 9.241569
Rin73_24 in73_23 in73_24 9.241569
Rin73_25 in73_24 in73_25 9.241569
Rin73_26 in73_25 in73_26 9.241569
Rin73_27 in73_26 in73_27 9.241569
Rin73_28 in73_27 in73_28 9.241569
Rin73_29 in73 in73_29 9.241569
Rin73_30 in73_29 in73_30 9.241569
Rin73_31 in73_30 in73_31 9.241569
Rin73_32 in73_31 in73_32 9.241569
Rin73_33 in73_32 in73_33 9.241569
Rin73_34 in73_33 in73_34 9.241569
Rin73_35 in73_34 in73_35 9.241569
Rin73_36 in73_35 in73_36 9.241569
Rin73_37 in73_36 in73_37 9.241569
Rin73_38 in73_37 in73_38 9.241569
Rin73_39 in73_38 in73_39 9.241569
Rin73_40 in73_39 in73_40 9.241569
Rin73_41 in73_40 in73_41 9.241569
Rin73_42 in73_41 in73_42 9.241569
Rin73_43 in73_42 in73_43 9.241569
Rin73_44 in73_43 in73_44 9.241569
Rin73_45 in73_44 in73_45 9.241569
Rin73_46 in73_45 in73_46 9.241569
Rin73_47 in73_46 in73_47 9.241569
Rin73_48 in73_47 in73_48 9.241569
Rin73_49 in73_48 in73_49 9.241569
Rin73_50 in73_49 in73_50 9.241569
Rin73_51 in73_50 in73_51 9.241569
Rin73_52 in73_51 in73_52 9.241569
Rin73_53 in73_52 in73_53 9.241569
Rin73_54 in73_53 in73_54 9.241569
Rin73_55 in73_54 in73_55 9.241569
Rin73_56 in73_55 in73_56 9.241569
Rin73_57 in73 in73_57 9.241569
Rin73_58 in73_57 in73_58 9.241569
Rin73_59 in73_58 in73_59 9.241569
Rin73_60 in73_59 in73_60 9.241569
Rin73_61 in73_60 in73_61 9.241569
Rin73_62 in73_61 in73_62 9.241569
Rin73_63 in73_62 in73_63 9.241569
Rin73_64 in73_63 in73_64 9.241569
Rin73_65 in73_64 in73_65 9.241569
Rin73_66 in73_65 in73_66 9.241569
Rin73_67 in73_66 in73_67 9.241569
Rin73_68 in73_67 in73_68 9.241569
Rin73_69 in73_68 in73_69 9.241569
Rin73_70 in73_69 in73_70 9.241569
Rin73_71 in73_70 in73_71 9.241569
Rin73_72 in73_71 in73_72 9.241569
Rin73_73 in73_72 in73_73 9.241569
Rin73_74 in73_73 in73_74 9.241569
Rin73_75 in73_74 in73_75 9.241569
Rin73_76 in73_75 in73_76 9.241569
Rin73_77 in73_76 in73_77 9.241569
Rin73_78 in73_77 in73_78 9.241569
Rin73_79 in73_78 in73_79 9.241569
Rin73_80 in73_79 in73_80 9.241569
Rin73_81 in73_80 in73_81 9.241569
Rin73_82 in73_81 in73_82 9.241569
Rin73_83 in73_82 in73_83 9.241569
Rin73_84 in73_83 in73_84 9.241569
Rin74_1 in74 in74_1 9.241569
Rin74_2 in74_1 in74_2 9.241569
Rin74_3 in74_2 in74_3 9.241569
Rin74_4 in74_3 in74_4 9.241569
Rin74_5 in74_4 in74_5 9.241569
Rin74_6 in74_5 in74_6 9.241569
Rin74_7 in74_6 in74_7 9.241569
Rin74_8 in74_7 in74_8 9.241569
Rin74_9 in74_8 in74_9 9.241569
Rin74_10 in74_9 in74_10 9.241569
Rin74_11 in74_10 in74_11 9.241569
Rin74_12 in74_11 in74_12 9.241569
Rin74_13 in74_12 in74_13 9.241569
Rin74_14 in74_13 in74_14 9.241569
Rin74_15 in74_14 in74_15 9.241569
Rin74_16 in74_15 in74_16 9.241569
Rin74_17 in74_16 in74_17 9.241569
Rin74_18 in74_17 in74_18 9.241569
Rin74_19 in74_18 in74_19 9.241569
Rin74_20 in74_19 in74_20 9.241569
Rin74_21 in74_20 in74_21 9.241569
Rin74_22 in74_21 in74_22 9.241569
Rin74_23 in74_22 in74_23 9.241569
Rin74_24 in74_23 in74_24 9.241569
Rin74_25 in74_24 in74_25 9.241569
Rin74_26 in74_25 in74_26 9.241569
Rin74_27 in74_26 in74_27 9.241569
Rin74_28 in74_27 in74_28 9.241569
Rin74_29 in74 in74_29 9.241569
Rin74_30 in74_29 in74_30 9.241569
Rin74_31 in74_30 in74_31 9.241569
Rin74_32 in74_31 in74_32 9.241569
Rin74_33 in74_32 in74_33 9.241569
Rin74_34 in74_33 in74_34 9.241569
Rin74_35 in74_34 in74_35 9.241569
Rin74_36 in74_35 in74_36 9.241569
Rin74_37 in74_36 in74_37 9.241569
Rin74_38 in74_37 in74_38 9.241569
Rin74_39 in74_38 in74_39 9.241569
Rin74_40 in74_39 in74_40 9.241569
Rin74_41 in74_40 in74_41 9.241569
Rin74_42 in74_41 in74_42 9.241569
Rin74_43 in74_42 in74_43 9.241569
Rin74_44 in74_43 in74_44 9.241569
Rin74_45 in74_44 in74_45 9.241569
Rin74_46 in74_45 in74_46 9.241569
Rin74_47 in74_46 in74_47 9.241569
Rin74_48 in74_47 in74_48 9.241569
Rin74_49 in74_48 in74_49 9.241569
Rin74_50 in74_49 in74_50 9.241569
Rin74_51 in74_50 in74_51 9.241569
Rin74_52 in74_51 in74_52 9.241569
Rin74_53 in74_52 in74_53 9.241569
Rin74_54 in74_53 in74_54 9.241569
Rin74_55 in74_54 in74_55 9.241569
Rin74_56 in74_55 in74_56 9.241569
Rin74_57 in74 in74_57 9.241569
Rin74_58 in74_57 in74_58 9.241569
Rin74_59 in74_58 in74_59 9.241569
Rin74_60 in74_59 in74_60 9.241569
Rin74_61 in74_60 in74_61 9.241569
Rin74_62 in74_61 in74_62 9.241569
Rin74_63 in74_62 in74_63 9.241569
Rin74_64 in74_63 in74_64 9.241569
Rin74_65 in74_64 in74_65 9.241569
Rin74_66 in74_65 in74_66 9.241569
Rin74_67 in74_66 in74_67 9.241569
Rin74_68 in74_67 in74_68 9.241569
Rin74_69 in74_68 in74_69 9.241569
Rin74_70 in74_69 in74_70 9.241569
Rin74_71 in74_70 in74_71 9.241569
Rin74_72 in74_71 in74_72 9.241569
Rin74_73 in74_72 in74_73 9.241569
Rin74_74 in74_73 in74_74 9.241569
Rin74_75 in74_74 in74_75 9.241569
Rin74_76 in74_75 in74_76 9.241569
Rin74_77 in74_76 in74_77 9.241569
Rin74_78 in74_77 in74_78 9.241569
Rin74_79 in74_78 in74_79 9.241569
Rin74_80 in74_79 in74_80 9.241569
Rin74_81 in74_80 in74_81 9.241569
Rin74_82 in74_81 in74_82 9.241569
Rin74_83 in74_82 in74_83 9.241569
Rin74_84 in74_83 in74_84 9.241569
Rin75_1 in75 in75_1 9.241569
Rin75_2 in75_1 in75_2 9.241569
Rin75_3 in75_2 in75_3 9.241569
Rin75_4 in75_3 in75_4 9.241569
Rin75_5 in75_4 in75_5 9.241569
Rin75_6 in75_5 in75_6 9.241569
Rin75_7 in75_6 in75_7 9.241569
Rin75_8 in75_7 in75_8 9.241569
Rin75_9 in75_8 in75_9 9.241569
Rin75_10 in75_9 in75_10 9.241569
Rin75_11 in75_10 in75_11 9.241569
Rin75_12 in75_11 in75_12 9.241569
Rin75_13 in75_12 in75_13 9.241569
Rin75_14 in75_13 in75_14 9.241569
Rin75_15 in75_14 in75_15 9.241569
Rin75_16 in75_15 in75_16 9.241569
Rin75_17 in75_16 in75_17 9.241569
Rin75_18 in75_17 in75_18 9.241569
Rin75_19 in75_18 in75_19 9.241569
Rin75_20 in75_19 in75_20 9.241569
Rin75_21 in75_20 in75_21 9.241569
Rin75_22 in75_21 in75_22 9.241569
Rin75_23 in75_22 in75_23 9.241569
Rin75_24 in75_23 in75_24 9.241569
Rin75_25 in75_24 in75_25 9.241569
Rin75_26 in75_25 in75_26 9.241569
Rin75_27 in75_26 in75_27 9.241569
Rin75_28 in75_27 in75_28 9.241569
Rin75_29 in75 in75_29 9.241569
Rin75_30 in75_29 in75_30 9.241569
Rin75_31 in75_30 in75_31 9.241569
Rin75_32 in75_31 in75_32 9.241569
Rin75_33 in75_32 in75_33 9.241569
Rin75_34 in75_33 in75_34 9.241569
Rin75_35 in75_34 in75_35 9.241569
Rin75_36 in75_35 in75_36 9.241569
Rin75_37 in75_36 in75_37 9.241569
Rin75_38 in75_37 in75_38 9.241569
Rin75_39 in75_38 in75_39 9.241569
Rin75_40 in75_39 in75_40 9.241569
Rin75_41 in75_40 in75_41 9.241569
Rin75_42 in75_41 in75_42 9.241569
Rin75_43 in75_42 in75_43 9.241569
Rin75_44 in75_43 in75_44 9.241569
Rin75_45 in75_44 in75_45 9.241569
Rin75_46 in75_45 in75_46 9.241569
Rin75_47 in75_46 in75_47 9.241569
Rin75_48 in75_47 in75_48 9.241569
Rin75_49 in75_48 in75_49 9.241569
Rin75_50 in75_49 in75_50 9.241569
Rin75_51 in75_50 in75_51 9.241569
Rin75_52 in75_51 in75_52 9.241569
Rin75_53 in75_52 in75_53 9.241569
Rin75_54 in75_53 in75_54 9.241569
Rin75_55 in75_54 in75_55 9.241569
Rin75_56 in75_55 in75_56 9.241569
Rin75_57 in75 in75_57 9.241569
Rin75_58 in75_57 in75_58 9.241569
Rin75_59 in75_58 in75_59 9.241569
Rin75_60 in75_59 in75_60 9.241569
Rin75_61 in75_60 in75_61 9.241569
Rin75_62 in75_61 in75_62 9.241569
Rin75_63 in75_62 in75_63 9.241569
Rin75_64 in75_63 in75_64 9.241569
Rin75_65 in75_64 in75_65 9.241569
Rin75_66 in75_65 in75_66 9.241569
Rin75_67 in75_66 in75_67 9.241569
Rin75_68 in75_67 in75_68 9.241569
Rin75_69 in75_68 in75_69 9.241569
Rin75_70 in75_69 in75_70 9.241569
Rin75_71 in75_70 in75_71 9.241569
Rin75_72 in75_71 in75_72 9.241569
Rin75_73 in75_72 in75_73 9.241569
Rin75_74 in75_73 in75_74 9.241569
Rin75_75 in75_74 in75_75 9.241569
Rin75_76 in75_75 in75_76 9.241569
Rin75_77 in75_76 in75_77 9.241569
Rin75_78 in75_77 in75_78 9.241569
Rin75_79 in75_78 in75_79 9.241569
Rin75_80 in75_79 in75_80 9.241569
Rin75_81 in75_80 in75_81 9.241569
Rin75_82 in75_81 in75_82 9.241569
Rin75_83 in75_82 in75_83 9.241569
Rin75_84 in75_83 in75_84 9.241569
Rin76_1 in76 in76_1 9.241569
Rin76_2 in76_1 in76_2 9.241569
Rin76_3 in76_2 in76_3 9.241569
Rin76_4 in76_3 in76_4 9.241569
Rin76_5 in76_4 in76_5 9.241569
Rin76_6 in76_5 in76_6 9.241569
Rin76_7 in76_6 in76_7 9.241569
Rin76_8 in76_7 in76_8 9.241569
Rin76_9 in76_8 in76_9 9.241569
Rin76_10 in76_9 in76_10 9.241569
Rin76_11 in76_10 in76_11 9.241569
Rin76_12 in76_11 in76_12 9.241569
Rin76_13 in76_12 in76_13 9.241569
Rin76_14 in76_13 in76_14 9.241569
Rin76_15 in76_14 in76_15 9.241569
Rin76_16 in76_15 in76_16 9.241569
Rin76_17 in76_16 in76_17 9.241569
Rin76_18 in76_17 in76_18 9.241569
Rin76_19 in76_18 in76_19 9.241569
Rin76_20 in76_19 in76_20 9.241569
Rin76_21 in76_20 in76_21 9.241569
Rin76_22 in76_21 in76_22 9.241569
Rin76_23 in76_22 in76_23 9.241569
Rin76_24 in76_23 in76_24 9.241569
Rin76_25 in76_24 in76_25 9.241569
Rin76_26 in76_25 in76_26 9.241569
Rin76_27 in76_26 in76_27 9.241569
Rin76_28 in76_27 in76_28 9.241569
Rin76_29 in76 in76_29 9.241569
Rin76_30 in76_29 in76_30 9.241569
Rin76_31 in76_30 in76_31 9.241569
Rin76_32 in76_31 in76_32 9.241569
Rin76_33 in76_32 in76_33 9.241569
Rin76_34 in76_33 in76_34 9.241569
Rin76_35 in76_34 in76_35 9.241569
Rin76_36 in76_35 in76_36 9.241569
Rin76_37 in76_36 in76_37 9.241569
Rin76_38 in76_37 in76_38 9.241569
Rin76_39 in76_38 in76_39 9.241569
Rin76_40 in76_39 in76_40 9.241569
Rin76_41 in76_40 in76_41 9.241569
Rin76_42 in76_41 in76_42 9.241569
Rin76_43 in76_42 in76_43 9.241569
Rin76_44 in76_43 in76_44 9.241569
Rin76_45 in76_44 in76_45 9.241569
Rin76_46 in76_45 in76_46 9.241569
Rin76_47 in76_46 in76_47 9.241569
Rin76_48 in76_47 in76_48 9.241569
Rin76_49 in76_48 in76_49 9.241569
Rin76_50 in76_49 in76_50 9.241569
Rin76_51 in76_50 in76_51 9.241569
Rin76_52 in76_51 in76_52 9.241569
Rin76_53 in76_52 in76_53 9.241569
Rin76_54 in76_53 in76_54 9.241569
Rin76_55 in76_54 in76_55 9.241569
Rin76_56 in76_55 in76_56 9.241569
Rin76_57 in76 in76_57 9.241569
Rin76_58 in76_57 in76_58 9.241569
Rin76_59 in76_58 in76_59 9.241569
Rin76_60 in76_59 in76_60 9.241569
Rin76_61 in76_60 in76_61 9.241569
Rin76_62 in76_61 in76_62 9.241569
Rin76_63 in76_62 in76_63 9.241569
Rin76_64 in76_63 in76_64 9.241569
Rin76_65 in76_64 in76_65 9.241569
Rin76_66 in76_65 in76_66 9.241569
Rin76_67 in76_66 in76_67 9.241569
Rin76_68 in76_67 in76_68 9.241569
Rin76_69 in76_68 in76_69 9.241569
Rin76_70 in76_69 in76_70 9.241569
Rin76_71 in76_70 in76_71 9.241569
Rin76_72 in76_71 in76_72 9.241569
Rin76_73 in76_72 in76_73 9.241569
Rin76_74 in76_73 in76_74 9.241569
Rin76_75 in76_74 in76_75 9.241569
Rin76_76 in76_75 in76_76 9.241569
Rin76_77 in76_76 in76_77 9.241569
Rin76_78 in76_77 in76_78 9.241569
Rin76_79 in76_78 in76_79 9.241569
Rin76_80 in76_79 in76_80 9.241569
Rin76_81 in76_80 in76_81 9.241569
Rin76_82 in76_81 in76_82 9.241569
Rin76_83 in76_82 in76_83 9.241569
Rin76_84 in76_83 in76_84 9.241569
Rin77_1 in77 in77_1 9.241569
Rin77_2 in77_1 in77_2 9.241569
Rin77_3 in77_2 in77_3 9.241569
Rin77_4 in77_3 in77_4 9.241569
Rin77_5 in77_4 in77_5 9.241569
Rin77_6 in77_5 in77_6 9.241569
Rin77_7 in77_6 in77_7 9.241569
Rin77_8 in77_7 in77_8 9.241569
Rin77_9 in77_8 in77_9 9.241569
Rin77_10 in77_9 in77_10 9.241569
Rin77_11 in77_10 in77_11 9.241569
Rin77_12 in77_11 in77_12 9.241569
Rin77_13 in77_12 in77_13 9.241569
Rin77_14 in77_13 in77_14 9.241569
Rin77_15 in77_14 in77_15 9.241569
Rin77_16 in77_15 in77_16 9.241569
Rin77_17 in77_16 in77_17 9.241569
Rin77_18 in77_17 in77_18 9.241569
Rin77_19 in77_18 in77_19 9.241569
Rin77_20 in77_19 in77_20 9.241569
Rin77_21 in77_20 in77_21 9.241569
Rin77_22 in77_21 in77_22 9.241569
Rin77_23 in77_22 in77_23 9.241569
Rin77_24 in77_23 in77_24 9.241569
Rin77_25 in77_24 in77_25 9.241569
Rin77_26 in77_25 in77_26 9.241569
Rin77_27 in77_26 in77_27 9.241569
Rin77_28 in77_27 in77_28 9.241569
Rin77_29 in77 in77_29 9.241569
Rin77_30 in77_29 in77_30 9.241569
Rin77_31 in77_30 in77_31 9.241569
Rin77_32 in77_31 in77_32 9.241569
Rin77_33 in77_32 in77_33 9.241569
Rin77_34 in77_33 in77_34 9.241569
Rin77_35 in77_34 in77_35 9.241569
Rin77_36 in77_35 in77_36 9.241569
Rin77_37 in77_36 in77_37 9.241569
Rin77_38 in77_37 in77_38 9.241569
Rin77_39 in77_38 in77_39 9.241569
Rin77_40 in77_39 in77_40 9.241569
Rin77_41 in77_40 in77_41 9.241569
Rin77_42 in77_41 in77_42 9.241569
Rin77_43 in77_42 in77_43 9.241569
Rin77_44 in77_43 in77_44 9.241569
Rin77_45 in77_44 in77_45 9.241569
Rin77_46 in77_45 in77_46 9.241569
Rin77_47 in77_46 in77_47 9.241569
Rin77_48 in77_47 in77_48 9.241569
Rin77_49 in77_48 in77_49 9.241569
Rin77_50 in77_49 in77_50 9.241569
Rin77_51 in77_50 in77_51 9.241569
Rin77_52 in77_51 in77_52 9.241569
Rin77_53 in77_52 in77_53 9.241569
Rin77_54 in77_53 in77_54 9.241569
Rin77_55 in77_54 in77_55 9.241569
Rin77_56 in77_55 in77_56 9.241569
Rin77_57 in77 in77_57 9.241569
Rin77_58 in77_57 in77_58 9.241569
Rin77_59 in77_58 in77_59 9.241569
Rin77_60 in77_59 in77_60 9.241569
Rin77_61 in77_60 in77_61 9.241569
Rin77_62 in77_61 in77_62 9.241569
Rin77_63 in77_62 in77_63 9.241569
Rin77_64 in77_63 in77_64 9.241569
Rin77_65 in77_64 in77_65 9.241569
Rin77_66 in77_65 in77_66 9.241569
Rin77_67 in77_66 in77_67 9.241569
Rin77_68 in77_67 in77_68 9.241569
Rin77_69 in77_68 in77_69 9.241569
Rin77_70 in77_69 in77_70 9.241569
Rin77_71 in77_70 in77_71 9.241569
Rin77_72 in77_71 in77_72 9.241569
Rin77_73 in77_72 in77_73 9.241569
Rin77_74 in77_73 in77_74 9.241569
Rin77_75 in77_74 in77_75 9.241569
Rin77_76 in77_75 in77_76 9.241569
Rin77_77 in77_76 in77_77 9.241569
Rin77_78 in77_77 in77_78 9.241569
Rin77_79 in77_78 in77_79 9.241569
Rin77_80 in77_79 in77_80 9.241569
Rin77_81 in77_80 in77_81 9.241569
Rin77_82 in77_81 in77_82 9.241569
Rin77_83 in77_82 in77_83 9.241569
Rin77_84 in77_83 in77_84 9.241569
Rin78_1 in78 in78_1 9.241569
Rin78_2 in78_1 in78_2 9.241569
Rin78_3 in78_2 in78_3 9.241569
Rin78_4 in78_3 in78_4 9.241569
Rin78_5 in78_4 in78_5 9.241569
Rin78_6 in78_5 in78_6 9.241569
Rin78_7 in78_6 in78_7 9.241569
Rin78_8 in78_7 in78_8 9.241569
Rin78_9 in78_8 in78_9 9.241569
Rin78_10 in78_9 in78_10 9.241569
Rin78_11 in78_10 in78_11 9.241569
Rin78_12 in78_11 in78_12 9.241569
Rin78_13 in78_12 in78_13 9.241569
Rin78_14 in78_13 in78_14 9.241569
Rin78_15 in78_14 in78_15 9.241569
Rin78_16 in78_15 in78_16 9.241569
Rin78_17 in78_16 in78_17 9.241569
Rin78_18 in78_17 in78_18 9.241569
Rin78_19 in78_18 in78_19 9.241569
Rin78_20 in78_19 in78_20 9.241569
Rin78_21 in78_20 in78_21 9.241569
Rin78_22 in78_21 in78_22 9.241569
Rin78_23 in78_22 in78_23 9.241569
Rin78_24 in78_23 in78_24 9.241569
Rin78_25 in78_24 in78_25 9.241569
Rin78_26 in78_25 in78_26 9.241569
Rin78_27 in78_26 in78_27 9.241569
Rin78_28 in78_27 in78_28 9.241569
Rin78_29 in78 in78_29 9.241569
Rin78_30 in78_29 in78_30 9.241569
Rin78_31 in78_30 in78_31 9.241569
Rin78_32 in78_31 in78_32 9.241569
Rin78_33 in78_32 in78_33 9.241569
Rin78_34 in78_33 in78_34 9.241569
Rin78_35 in78_34 in78_35 9.241569
Rin78_36 in78_35 in78_36 9.241569
Rin78_37 in78_36 in78_37 9.241569
Rin78_38 in78_37 in78_38 9.241569
Rin78_39 in78_38 in78_39 9.241569
Rin78_40 in78_39 in78_40 9.241569
Rin78_41 in78_40 in78_41 9.241569
Rin78_42 in78_41 in78_42 9.241569
Rin78_43 in78_42 in78_43 9.241569
Rin78_44 in78_43 in78_44 9.241569
Rin78_45 in78_44 in78_45 9.241569
Rin78_46 in78_45 in78_46 9.241569
Rin78_47 in78_46 in78_47 9.241569
Rin78_48 in78_47 in78_48 9.241569
Rin78_49 in78_48 in78_49 9.241569
Rin78_50 in78_49 in78_50 9.241569
Rin78_51 in78_50 in78_51 9.241569
Rin78_52 in78_51 in78_52 9.241569
Rin78_53 in78_52 in78_53 9.241569
Rin78_54 in78_53 in78_54 9.241569
Rin78_55 in78_54 in78_55 9.241569
Rin78_56 in78_55 in78_56 9.241569
Rin78_57 in78 in78_57 9.241569
Rin78_58 in78_57 in78_58 9.241569
Rin78_59 in78_58 in78_59 9.241569
Rin78_60 in78_59 in78_60 9.241569
Rin78_61 in78_60 in78_61 9.241569
Rin78_62 in78_61 in78_62 9.241569
Rin78_63 in78_62 in78_63 9.241569
Rin78_64 in78_63 in78_64 9.241569
Rin78_65 in78_64 in78_65 9.241569
Rin78_66 in78_65 in78_66 9.241569
Rin78_67 in78_66 in78_67 9.241569
Rin78_68 in78_67 in78_68 9.241569
Rin78_69 in78_68 in78_69 9.241569
Rin78_70 in78_69 in78_70 9.241569
Rin78_71 in78_70 in78_71 9.241569
Rin78_72 in78_71 in78_72 9.241569
Rin78_73 in78_72 in78_73 9.241569
Rin78_74 in78_73 in78_74 9.241569
Rin78_75 in78_74 in78_75 9.241569
Rin78_76 in78_75 in78_76 9.241569
Rin78_77 in78_76 in78_77 9.241569
Rin78_78 in78_77 in78_78 9.241569
Rin78_79 in78_78 in78_79 9.241569
Rin78_80 in78_79 in78_80 9.241569
Rin78_81 in78_80 in78_81 9.241569
Rin78_82 in78_81 in78_82 9.241569
Rin78_83 in78_82 in78_83 9.241569
Rin78_84 in78_83 in78_84 9.241569
Rin79_1 in79 in79_1 9.241569
Rin79_2 in79_1 in79_2 9.241569
Rin79_3 in79_2 in79_3 9.241569
Rin79_4 in79_3 in79_4 9.241569
Rin79_5 in79_4 in79_5 9.241569
Rin79_6 in79_5 in79_6 9.241569
Rin79_7 in79_6 in79_7 9.241569
Rin79_8 in79_7 in79_8 9.241569
Rin79_9 in79_8 in79_9 9.241569
Rin79_10 in79_9 in79_10 9.241569
Rin79_11 in79_10 in79_11 9.241569
Rin79_12 in79_11 in79_12 9.241569
Rin79_13 in79_12 in79_13 9.241569
Rin79_14 in79_13 in79_14 9.241569
Rin79_15 in79_14 in79_15 9.241569
Rin79_16 in79_15 in79_16 9.241569
Rin79_17 in79_16 in79_17 9.241569
Rin79_18 in79_17 in79_18 9.241569
Rin79_19 in79_18 in79_19 9.241569
Rin79_20 in79_19 in79_20 9.241569
Rin79_21 in79_20 in79_21 9.241569
Rin79_22 in79_21 in79_22 9.241569
Rin79_23 in79_22 in79_23 9.241569
Rin79_24 in79_23 in79_24 9.241569
Rin79_25 in79_24 in79_25 9.241569
Rin79_26 in79_25 in79_26 9.241569
Rin79_27 in79_26 in79_27 9.241569
Rin79_28 in79_27 in79_28 9.241569
Rin79_29 in79 in79_29 9.241569
Rin79_30 in79_29 in79_30 9.241569
Rin79_31 in79_30 in79_31 9.241569
Rin79_32 in79_31 in79_32 9.241569
Rin79_33 in79_32 in79_33 9.241569
Rin79_34 in79_33 in79_34 9.241569
Rin79_35 in79_34 in79_35 9.241569
Rin79_36 in79_35 in79_36 9.241569
Rin79_37 in79_36 in79_37 9.241569
Rin79_38 in79_37 in79_38 9.241569
Rin79_39 in79_38 in79_39 9.241569
Rin79_40 in79_39 in79_40 9.241569
Rin79_41 in79_40 in79_41 9.241569
Rin79_42 in79_41 in79_42 9.241569
Rin79_43 in79_42 in79_43 9.241569
Rin79_44 in79_43 in79_44 9.241569
Rin79_45 in79_44 in79_45 9.241569
Rin79_46 in79_45 in79_46 9.241569
Rin79_47 in79_46 in79_47 9.241569
Rin79_48 in79_47 in79_48 9.241569
Rin79_49 in79_48 in79_49 9.241569
Rin79_50 in79_49 in79_50 9.241569
Rin79_51 in79_50 in79_51 9.241569
Rin79_52 in79_51 in79_52 9.241569
Rin79_53 in79_52 in79_53 9.241569
Rin79_54 in79_53 in79_54 9.241569
Rin79_55 in79_54 in79_55 9.241569
Rin79_56 in79_55 in79_56 9.241569
Rin79_57 in79 in79_57 9.241569
Rin79_58 in79_57 in79_58 9.241569
Rin79_59 in79_58 in79_59 9.241569
Rin79_60 in79_59 in79_60 9.241569
Rin79_61 in79_60 in79_61 9.241569
Rin79_62 in79_61 in79_62 9.241569
Rin79_63 in79_62 in79_63 9.241569
Rin79_64 in79_63 in79_64 9.241569
Rin79_65 in79_64 in79_65 9.241569
Rin79_66 in79_65 in79_66 9.241569
Rin79_67 in79_66 in79_67 9.241569
Rin79_68 in79_67 in79_68 9.241569
Rin79_69 in79_68 in79_69 9.241569
Rin79_70 in79_69 in79_70 9.241569
Rin79_71 in79_70 in79_71 9.241569
Rin79_72 in79_71 in79_72 9.241569
Rin79_73 in79_72 in79_73 9.241569
Rin79_74 in79_73 in79_74 9.241569
Rin79_75 in79_74 in79_75 9.241569
Rin79_76 in79_75 in79_76 9.241569
Rin79_77 in79_76 in79_77 9.241569
Rin79_78 in79_77 in79_78 9.241569
Rin79_79 in79_78 in79_79 9.241569
Rin79_80 in79_79 in79_80 9.241569
Rin79_81 in79_80 in79_81 9.241569
Rin79_82 in79_81 in79_82 9.241569
Rin79_83 in79_82 in79_83 9.241569
Rin79_84 in79_83 in79_84 9.241569
Rin80_1 in80 in80_1 9.241569
Rin80_2 in80_1 in80_2 9.241569
Rin80_3 in80_2 in80_3 9.241569
Rin80_4 in80_3 in80_4 9.241569
Rin80_5 in80_4 in80_5 9.241569
Rin80_6 in80_5 in80_6 9.241569
Rin80_7 in80_6 in80_7 9.241569
Rin80_8 in80_7 in80_8 9.241569
Rin80_9 in80_8 in80_9 9.241569
Rin80_10 in80_9 in80_10 9.241569
Rin80_11 in80_10 in80_11 9.241569
Rin80_12 in80_11 in80_12 9.241569
Rin80_13 in80_12 in80_13 9.241569
Rin80_14 in80_13 in80_14 9.241569
Rin80_15 in80_14 in80_15 9.241569
Rin80_16 in80_15 in80_16 9.241569
Rin80_17 in80_16 in80_17 9.241569
Rin80_18 in80_17 in80_18 9.241569
Rin80_19 in80_18 in80_19 9.241569
Rin80_20 in80_19 in80_20 9.241569
Rin80_21 in80_20 in80_21 9.241569
Rin80_22 in80_21 in80_22 9.241569
Rin80_23 in80_22 in80_23 9.241569
Rin80_24 in80_23 in80_24 9.241569
Rin80_25 in80_24 in80_25 9.241569
Rin80_26 in80_25 in80_26 9.241569
Rin80_27 in80_26 in80_27 9.241569
Rin80_28 in80_27 in80_28 9.241569
Rin80_29 in80 in80_29 9.241569
Rin80_30 in80_29 in80_30 9.241569
Rin80_31 in80_30 in80_31 9.241569
Rin80_32 in80_31 in80_32 9.241569
Rin80_33 in80_32 in80_33 9.241569
Rin80_34 in80_33 in80_34 9.241569
Rin80_35 in80_34 in80_35 9.241569
Rin80_36 in80_35 in80_36 9.241569
Rin80_37 in80_36 in80_37 9.241569
Rin80_38 in80_37 in80_38 9.241569
Rin80_39 in80_38 in80_39 9.241569
Rin80_40 in80_39 in80_40 9.241569
Rin80_41 in80_40 in80_41 9.241569
Rin80_42 in80_41 in80_42 9.241569
Rin80_43 in80_42 in80_43 9.241569
Rin80_44 in80_43 in80_44 9.241569
Rin80_45 in80_44 in80_45 9.241569
Rin80_46 in80_45 in80_46 9.241569
Rin80_47 in80_46 in80_47 9.241569
Rin80_48 in80_47 in80_48 9.241569
Rin80_49 in80_48 in80_49 9.241569
Rin80_50 in80_49 in80_50 9.241569
Rin80_51 in80_50 in80_51 9.241569
Rin80_52 in80_51 in80_52 9.241569
Rin80_53 in80_52 in80_53 9.241569
Rin80_54 in80_53 in80_54 9.241569
Rin80_55 in80_54 in80_55 9.241569
Rin80_56 in80_55 in80_56 9.241569
Rin80_57 in80 in80_57 9.241569
Rin80_58 in80_57 in80_58 9.241569
Rin80_59 in80_58 in80_59 9.241569
Rin80_60 in80_59 in80_60 9.241569
Rin80_61 in80_60 in80_61 9.241569
Rin80_62 in80_61 in80_62 9.241569
Rin80_63 in80_62 in80_63 9.241569
Rin80_64 in80_63 in80_64 9.241569
Rin80_65 in80_64 in80_65 9.241569
Rin80_66 in80_65 in80_66 9.241569
Rin80_67 in80_66 in80_67 9.241569
Rin80_68 in80_67 in80_68 9.241569
Rin80_69 in80_68 in80_69 9.241569
Rin80_70 in80_69 in80_70 9.241569
Rin80_71 in80_70 in80_71 9.241569
Rin80_72 in80_71 in80_72 9.241569
Rin80_73 in80_72 in80_73 9.241569
Rin80_74 in80_73 in80_74 9.241569
Rin80_75 in80_74 in80_75 9.241569
Rin80_76 in80_75 in80_76 9.241569
Rin80_77 in80_76 in80_77 9.241569
Rin80_78 in80_77 in80_78 9.241569
Rin80_79 in80_78 in80_79 9.241569
Rin80_80 in80_79 in80_80 9.241569
Rin80_81 in80_80 in80_81 9.241569
Rin80_82 in80_81 in80_82 9.241569
Rin80_83 in80_82 in80_83 9.241569
Rin80_84 in80_83 in80_84 9.241569
Rin81_1 in81 in81_1 9.241569
Rin81_2 in81_1 in81_2 9.241569
Rin81_3 in81_2 in81_3 9.241569
Rin81_4 in81_3 in81_4 9.241569
Rin81_5 in81_4 in81_5 9.241569
Rin81_6 in81_5 in81_6 9.241569
Rin81_7 in81_6 in81_7 9.241569
Rin81_8 in81_7 in81_8 9.241569
Rin81_9 in81_8 in81_9 9.241569
Rin81_10 in81_9 in81_10 9.241569
Rin81_11 in81_10 in81_11 9.241569
Rin81_12 in81_11 in81_12 9.241569
Rin81_13 in81_12 in81_13 9.241569
Rin81_14 in81_13 in81_14 9.241569
Rin81_15 in81_14 in81_15 9.241569
Rin81_16 in81_15 in81_16 9.241569
Rin81_17 in81_16 in81_17 9.241569
Rin81_18 in81_17 in81_18 9.241569
Rin81_19 in81_18 in81_19 9.241569
Rin81_20 in81_19 in81_20 9.241569
Rin81_21 in81_20 in81_21 9.241569
Rin81_22 in81_21 in81_22 9.241569
Rin81_23 in81_22 in81_23 9.241569
Rin81_24 in81_23 in81_24 9.241569
Rin81_25 in81_24 in81_25 9.241569
Rin81_26 in81_25 in81_26 9.241569
Rin81_27 in81_26 in81_27 9.241569
Rin81_28 in81_27 in81_28 9.241569
Rin81_29 in81 in81_29 9.241569
Rin81_30 in81_29 in81_30 9.241569
Rin81_31 in81_30 in81_31 9.241569
Rin81_32 in81_31 in81_32 9.241569
Rin81_33 in81_32 in81_33 9.241569
Rin81_34 in81_33 in81_34 9.241569
Rin81_35 in81_34 in81_35 9.241569
Rin81_36 in81_35 in81_36 9.241569
Rin81_37 in81_36 in81_37 9.241569
Rin81_38 in81_37 in81_38 9.241569
Rin81_39 in81_38 in81_39 9.241569
Rin81_40 in81_39 in81_40 9.241569
Rin81_41 in81_40 in81_41 9.241569
Rin81_42 in81_41 in81_42 9.241569
Rin81_43 in81_42 in81_43 9.241569
Rin81_44 in81_43 in81_44 9.241569
Rin81_45 in81_44 in81_45 9.241569
Rin81_46 in81_45 in81_46 9.241569
Rin81_47 in81_46 in81_47 9.241569
Rin81_48 in81_47 in81_48 9.241569
Rin81_49 in81_48 in81_49 9.241569
Rin81_50 in81_49 in81_50 9.241569
Rin81_51 in81_50 in81_51 9.241569
Rin81_52 in81_51 in81_52 9.241569
Rin81_53 in81_52 in81_53 9.241569
Rin81_54 in81_53 in81_54 9.241569
Rin81_55 in81_54 in81_55 9.241569
Rin81_56 in81_55 in81_56 9.241569
Rin81_57 in81 in81_57 9.241569
Rin81_58 in81_57 in81_58 9.241569
Rin81_59 in81_58 in81_59 9.241569
Rin81_60 in81_59 in81_60 9.241569
Rin81_61 in81_60 in81_61 9.241569
Rin81_62 in81_61 in81_62 9.241569
Rin81_63 in81_62 in81_63 9.241569
Rin81_64 in81_63 in81_64 9.241569
Rin81_65 in81_64 in81_65 9.241569
Rin81_66 in81_65 in81_66 9.241569
Rin81_67 in81_66 in81_67 9.241569
Rin81_68 in81_67 in81_68 9.241569
Rin81_69 in81_68 in81_69 9.241569
Rin81_70 in81_69 in81_70 9.241569
Rin81_71 in81_70 in81_71 9.241569
Rin81_72 in81_71 in81_72 9.241569
Rin81_73 in81_72 in81_73 9.241569
Rin81_74 in81_73 in81_74 9.241569
Rin81_75 in81_74 in81_75 9.241569
Rin81_76 in81_75 in81_76 9.241569
Rin81_77 in81_76 in81_77 9.241569
Rin81_78 in81_77 in81_78 9.241569
Rin81_79 in81_78 in81_79 9.241569
Rin81_80 in81_79 in81_80 9.241569
Rin81_81 in81_80 in81_81 9.241569
Rin81_82 in81_81 in81_82 9.241569
Rin81_83 in81_82 in81_83 9.241569
Rin81_84 in81_83 in81_84 9.241569
Rin82_1 in82 in82_1 9.241569
Rin82_2 in82_1 in82_2 9.241569
Rin82_3 in82_2 in82_3 9.241569
Rin82_4 in82_3 in82_4 9.241569
Rin82_5 in82_4 in82_5 9.241569
Rin82_6 in82_5 in82_6 9.241569
Rin82_7 in82_6 in82_7 9.241569
Rin82_8 in82_7 in82_8 9.241569
Rin82_9 in82_8 in82_9 9.241569
Rin82_10 in82_9 in82_10 9.241569
Rin82_11 in82_10 in82_11 9.241569
Rin82_12 in82_11 in82_12 9.241569
Rin82_13 in82_12 in82_13 9.241569
Rin82_14 in82_13 in82_14 9.241569
Rin82_15 in82_14 in82_15 9.241569
Rin82_16 in82_15 in82_16 9.241569
Rin82_17 in82_16 in82_17 9.241569
Rin82_18 in82_17 in82_18 9.241569
Rin82_19 in82_18 in82_19 9.241569
Rin82_20 in82_19 in82_20 9.241569
Rin82_21 in82_20 in82_21 9.241569
Rin82_22 in82_21 in82_22 9.241569
Rin82_23 in82_22 in82_23 9.241569
Rin82_24 in82_23 in82_24 9.241569
Rin82_25 in82_24 in82_25 9.241569
Rin82_26 in82_25 in82_26 9.241569
Rin82_27 in82_26 in82_27 9.241569
Rin82_28 in82_27 in82_28 9.241569
Rin82_29 in82 in82_29 9.241569
Rin82_30 in82_29 in82_30 9.241569
Rin82_31 in82_30 in82_31 9.241569
Rin82_32 in82_31 in82_32 9.241569
Rin82_33 in82_32 in82_33 9.241569
Rin82_34 in82_33 in82_34 9.241569
Rin82_35 in82_34 in82_35 9.241569
Rin82_36 in82_35 in82_36 9.241569
Rin82_37 in82_36 in82_37 9.241569
Rin82_38 in82_37 in82_38 9.241569
Rin82_39 in82_38 in82_39 9.241569
Rin82_40 in82_39 in82_40 9.241569
Rin82_41 in82_40 in82_41 9.241569
Rin82_42 in82_41 in82_42 9.241569
Rin82_43 in82_42 in82_43 9.241569
Rin82_44 in82_43 in82_44 9.241569
Rin82_45 in82_44 in82_45 9.241569
Rin82_46 in82_45 in82_46 9.241569
Rin82_47 in82_46 in82_47 9.241569
Rin82_48 in82_47 in82_48 9.241569
Rin82_49 in82_48 in82_49 9.241569
Rin82_50 in82_49 in82_50 9.241569
Rin82_51 in82_50 in82_51 9.241569
Rin82_52 in82_51 in82_52 9.241569
Rin82_53 in82_52 in82_53 9.241569
Rin82_54 in82_53 in82_54 9.241569
Rin82_55 in82_54 in82_55 9.241569
Rin82_56 in82_55 in82_56 9.241569
Rin82_57 in82 in82_57 9.241569
Rin82_58 in82_57 in82_58 9.241569
Rin82_59 in82_58 in82_59 9.241569
Rin82_60 in82_59 in82_60 9.241569
Rin82_61 in82_60 in82_61 9.241569
Rin82_62 in82_61 in82_62 9.241569
Rin82_63 in82_62 in82_63 9.241569
Rin82_64 in82_63 in82_64 9.241569
Rin82_65 in82_64 in82_65 9.241569
Rin82_66 in82_65 in82_66 9.241569
Rin82_67 in82_66 in82_67 9.241569
Rin82_68 in82_67 in82_68 9.241569
Rin82_69 in82_68 in82_69 9.241569
Rin82_70 in82_69 in82_70 9.241569
Rin82_71 in82_70 in82_71 9.241569
Rin82_72 in82_71 in82_72 9.241569
Rin82_73 in82_72 in82_73 9.241569
Rin82_74 in82_73 in82_74 9.241569
Rin82_75 in82_74 in82_75 9.241569
Rin82_76 in82_75 in82_76 9.241569
Rin82_77 in82_76 in82_77 9.241569
Rin82_78 in82_77 in82_78 9.241569
Rin82_79 in82_78 in82_79 9.241569
Rin82_80 in82_79 in82_80 9.241569
Rin82_81 in82_80 in82_81 9.241569
Rin82_82 in82_81 in82_82 9.241569
Rin82_83 in82_82 in82_83 9.241569
Rin82_84 in82_83 in82_84 9.241569
Rin83_1 in83 in83_1 9.241569
Rin83_2 in83_1 in83_2 9.241569
Rin83_3 in83_2 in83_3 9.241569
Rin83_4 in83_3 in83_4 9.241569
Rin83_5 in83_4 in83_5 9.241569
Rin83_6 in83_5 in83_6 9.241569
Rin83_7 in83_6 in83_7 9.241569
Rin83_8 in83_7 in83_8 9.241569
Rin83_9 in83_8 in83_9 9.241569
Rin83_10 in83_9 in83_10 9.241569
Rin83_11 in83_10 in83_11 9.241569
Rin83_12 in83_11 in83_12 9.241569
Rin83_13 in83_12 in83_13 9.241569
Rin83_14 in83_13 in83_14 9.241569
Rin83_15 in83_14 in83_15 9.241569
Rin83_16 in83_15 in83_16 9.241569
Rin83_17 in83_16 in83_17 9.241569
Rin83_18 in83_17 in83_18 9.241569
Rin83_19 in83_18 in83_19 9.241569
Rin83_20 in83_19 in83_20 9.241569
Rin83_21 in83_20 in83_21 9.241569
Rin83_22 in83_21 in83_22 9.241569
Rin83_23 in83_22 in83_23 9.241569
Rin83_24 in83_23 in83_24 9.241569
Rin83_25 in83_24 in83_25 9.241569
Rin83_26 in83_25 in83_26 9.241569
Rin83_27 in83_26 in83_27 9.241569
Rin83_28 in83_27 in83_28 9.241569
Rin83_29 in83 in83_29 9.241569
Rin83_30 in83_29 in83_30 9.241569
Rin83_31 in83_30 in83_31 9.241569
Rin83_32 in83_31 in83_32 9.241569
Rin83_33 in83_32 in83_33 9.241569
Rin83_34 in83_33 in83_34 9.241569
Rin83_35 in83_34 in83_35 9.241569
Rin83_36 in83_35 in83_36 9.241569
Rin83_37 in83_36 in83_37 9.241569
Rin83_38 in83_37 in83_38 9.241569
Rin83_39 in83_38 in83_39 9.241569
Rin83_40 in83_39 in83_40 9.241569
Rin83_41 in83_40 in83_41 9.241569
Rin83_42 in83_41 in83_42 9.241569
Rin83_43 in83_42 in83_43 9.241569
Rin83_44 in83_43 in83_44 9.241569
Rin83_45 in83_44 in83_45 9.241569
Rin83_46 in83_45 in83_46 9.241569
Rin83_47 in83_46 in83_47 9.241569
Rin83_48 in83_47 in83_48 9.241569
Rin83_49 in83_48 in83_49 9.241569
Rin83_50 in83_49 in83_50 9.241569
Rin83_51 in83_50 in83_51 9.241569
Rin83_52 in83_51 in83_52 9.241569
Rin83_53 in83_52 in83_53 9.241569
Rin83_54 in83_53 in83_54 9.241569
Rin83_55 in83_54 in83_55 9.241569
Rin83_56 in83_55 in83_56 9.241569
Rin83_57 in83 in83_57 9.241569
Rin83_58 in83_57 in83_58 9.241569
Rin83_59 in83_58 in83_59 9.241569
Rin83_60 in83_59 in83_60 9.241569
Rin83_61 in83_60 in83_61 9.241569
Rin83_62 in83_61 in83_62 9.241569
Rin83_63 in83_62 in83_63 9.241569
Rin83_64 in83_63 in83_64 9.241569
Rin83_65 in83_64 in83_65 9.241569
Rin83_66 in83_65 in83_66 9.241569
Rin83_67 in83_66 in83_67 9.241569
Rin83_68 in83_67 in83_68 9.241569
Rin83_69 in83_68 in83_69 9.241569
Rin83_70 in83_69 in83_70 9.241569
Rin83_71 in83_70 in83_71 9.241569
Rin83_72 in83_71 in83_72 9.241569
Rin83_73 in83_72 in83_73 9.241569
Rin83_74 in83_73 in83_74 9.241569
Rin83_75 in83_74 in83_75 9.241569
Rin83_76 in83_75 in83_76 9.241569
Rin83_77 in83_76 in83_77 9.241569
Rin83_78 in83_77 in83_78 9.241569
Rin83_79 in83_78 in83_79 9.241569
Rin83_80 in83_79 in83_80 9.241569
Rin83_81 in83_80 in83_81 9.241569
Rin83_82 in83_81 in83_82 9.241569
Rin83_83 in83_82 in83_83 9.241569
Rin83_84 in83_83 in83_84 9.241569
Rin84_1 in84 in84_1 9.241569
Rin84_2 in84_1 in84_2 9.241569
Rin84_3 in84_2 in84_3 9.241569
Rin84_4 in84_3 in84_4 9.241569
Rin84_5 in84_4 in84_5 9.241569
Rin84_6 in84_5 in84_6 9.241569
Rin84_7 in84_6 in84_7 9.241569
Rin84_8 in84_7 in84_8 9.241569
Rin84_9 in84_8 in84_9 9.241569
Rin84_10 in84_9 in84_10 9.241569
Rin84_11 in84_10 in84_11 9.241569
Rin84_12 in84_11 in84_12 9.241569
Rin84_13 in84_12 in84_13 9.241569
Rin84_14 in84_13 in84_14 9.241569
Rin84_15 in84_14 in84_15 9.241569
Rin84_16 in84_15 in84_16 9.241569
Rin84_17 in84_16 in84_17 9.241569
Rin84_18 in84_17 in84_18 9.241569
Rin84_19 in84_18 in84_19 9.241569
Rin84_20 in84_19 in84_20 9.241569
Rin84_21 in84_20 in84_21 9.241569
Rin84_22 in84_21 in84_22 9.241569
Rin84_23 in84_22 in84_23 9.241569
Rin84_24 in84_23 in84_24 9.241569
Rin84_25 in84_24 in84_25 9.241569
Rin84_26 in84_25 in84_26 9.241569
Rin84_27 in84_26 in84_27 9.241569
Rin84_28 in84_27 in84_28 9.241569
Rin84_29 in84 in84_29 9.241569
Rin84_30 in84_29 in84_30 9.241569
Rin84_31 in84_30 in84_31 9.241569
Rin84_32 in84_31 in84_32 9.241569
Rin84_33 in84_32 in84_33 9.241569
Rin84_34 in84_33 in84_34 9.241569
Rin84_35 in84_34 in84_35 9.241569
Rin84_36 in84_35 in84_36 9.241569
Rin84_37 in84_36 in84_37 9.241569
Rin84_38 in84_37 in84_38 9.241569
Rin84_39 in84_38 in84_39 9.241569
Rin84_40 in84_39 in84_40 9.241569
Rin84_41 in84_40 in84_41 9.241569
Rin84_42 in84_41 in84_42 9.241569
Rin84_43 in84_42 in84_43 9.241569
Rin84_44 in84_43 in84_44 9.241569
Rin84_45 in84_44 in84_45 9.241569
Rin84_46 in84_45 in84_46 9.241569
Rin84_47 in84_46 in84_47 9.241569
Rin84_48 in84_47 in84_48 9.241569
Rin84_49 in84_48 in84_49 9.241569
Rin84_50 in84_49 in84_50 9.241569
Rin84_51 in84_50 in84_51 9.241569
Rin84_52 in84_51 in84_52 9.241569
Rin84_53 in84_52 in84_53 9.241569
Rin84_54 in84_53 in84_54 9.241569
Rin84_55 in84_54 in84_55 9.241569
Rin84_56 in84_55 in84_56 9.241569
Rin84_57 in84 in84_57 9.241569
Rin84_58 in84_57 in84_58 9.241569
Rin84_59 in84_58 in84_59 9.241569
Rin84_60 in84_59 in84_60 9.241569
Rin84_61 in84_60 in84_61 9.241569
Rin84_62 in84_61 in84_62 9.241569
Rin84_63 in84_62 in84_63 9.241569
Rin84_64 in84_63 in84_64 9.241569
Rin84_65 in84_64 in84_65 9.241569
Rin84_66 in84_65 in84_66 9.241569
Rin84_67 in84_66 in84_67 9.241569
Rin84_68 in84_67 in84_68 9.241569
Rin84_69 in84_68 in84_69 9.241569
Rin84_70 in84_69 in84_70 9.241569
Rin84_71 in84_70 in84_71 9.241569
Rin84_72 in84_71 in84_72 9.241569
Rin84_73 in84_72 in84_73 9.241569
Rin84_74 in84_73 in84_74 9.241569
Rin84_75 in84_74 in84_75 9.241569
Rin84_76 in84_75 in84_76 9.241569
Rin84_77 in84_76 in84_77 9.241569
Rin84_78 in84_77 in84_78 9.241569
Rin84_79 in84_78 in84_79 9.241569
Rin84_80 in84_79 in84_80 9.241569
Rin84_81 in84_80 in84_81 9.241569
Rin84_82 in84_81 in84_82 9.241569
Rin84_83 in84_82 in84_83 9.241569
Rin84_84 in84_83 in84_84 9.241569
Rin85_1 in85 in85_1 9.241569
Rin85_2 in85_1 in85_2 9.241569
Rin85_3 in85_2 in85_3 9.241569
Rin85_4 in85_3 in85_4 9.241569
Rin85_5 in85_4 in85_5 9.241569
Rin85_6 in85_5 in85_6 9.241569
Rin85_7 in85_6 in85_7 9.241569
Rin85_8 in85_7 in85_8 9.241569
Rin85_9 in85_8 in85_9 9.241569
Rin85_10 in85_9 in85_10 9.241569
Rin85_11 in85_10 in85_11 9.241569
Rin85_12 in85_11 in85_12 9.241569
Rin85_13 in85_12 in85_13 9.241569
Rin85_14 in85_13 in85_14 9.241569
Rin85_15 in85_14 in85_15 9.241569
Rin85_16 in85_15 in85_16 9.241569
Rin85_17 in85_16 in85_17 9.241569
Rin85_18 in85_17 in85_18 9.241569
Rin85_19 in85_18 in85_19 9.241569
Rin85_20 in85_19 in85_20 9.241569
Rin85_21 in85_20 in85_21 9.241569
Rin85_22 in85_21 in85_22 9.241569
Rin85_23 in85_22 in85_23 9.241569
Rin85_24 in85_23 in85_24 9.241569
Rin85_25 in85_24 in85_25 9.241569
Rin85_26 in85_25 in85_26 9.241569
Rin85_27 in85_26 in85_27 9.241569
Rin85_28 in85_27 in85_28 9.241569
Rin85_29 in85 in85_29 9.241569
Rin85_30 in85_29 in85_30 9.241569
Rin85_31 in85_30 in85_31 9.241569
Rin85_32 in85_31 in85_32 9.241569
Rin85_33 in85_32 in85_33 9.241569
Rin85_34 in85_33 in85_34 9.241569
Rin85_35 in85_34 in85_35 9.241569
Rin85_36 in85_35 in85_36 9.241569
Rin85_37 in85_36 in85_37 9.241569
Rin85_38 in85_37 in85_38 9.241569
Rin85_39 in85_38 in85_39 9.241569
Rin85_40 in85_39 in85_40 9.241569
Rin85_41 in85_40 in85_41 9.241569
Rin85_42 in85_41 in85_42 9.241569
Rin85_43 in85_42 in85_43 9.241569
Rin85_44 in85_43 in85_44 9.241569
Rin85_45 in85_44 in85_45 9.241569
Rin85_46 in85_45 in85_46 9.241569
Rin85_47 in85_46 in85_47 9.241569
Rin85_48 in85_47 in85_48 9.241569
Rin85_49 in85_48 in85_49 9.241569
Rin85_50 in85_49 in85_50 9.241569
Rin85_51 in85_50 in85_51 9.241569
Rin85_52 in85_51 in85_52 9.241569
Rin85_53 in85_52 in85_53 9.241569
Rin85_54 in85_53 in85_54 9.241569
Rin85_55 in85_54 in85_55 9.241569
Rin85_56 in85_55 in85_56 9.241569
Rin85_57 in85 in85_57 9.241569
Rin85_58 in85_57 in85_58 9.241569
Rin85_59 in85_58 in85_59 9.241569
Rin85_60 in85_59 in85_60 9.241569
Rin85_61 in85_60 in85_61 9.241569
Rin85_62 in85_61 in85_62 9.241569
Rin85_63 in85_62 in85_63 9.241569
Rin85_64 in85_63 in85_64 9.241569
Rin85_65 in85_64 in85_65 9.241569
Rin85_66 in85_65 in85_66 9.241569
Rin85_67 in85_66 in85_67 9.241569
Rin85_68 in85_67 in85_68 9.241569
Rin85_69 in85_68 in85_69 9.241569
Rin85_70 in85_69 in85_70 9.241569
Rin85_71 in85_70 in85_71 9.241569
Rin85_72 in85_71 in85_72 9.241569
Rin85_73 in85_72 in85_73 9.241569
Rin85_74 in85_73 in85_74 9.241569
Rin85_75 in85_74 in85_75 9.241569
Rin85_76 in85_75 in85_76 9.241569
Rin85_77 in85_76 in85_77 9.241569
Rin85_78 in85_77 in85_78 9.241569
Rin85_79 in85_78 in85_79 9.241569
Rin85_80 in85_79 in85_80 9.241569
Rin85_81 in85_80 in85_81 9.241569
Rin85_82 in85_81 in85_82 9.241569
Rin85_83 in85_82 in85_83 9.241569
Rin85_84 in85_83 in85_84 9.241569
Rin86_1 in86 in86_1 9.241569
Rin86_2 in86_1 in86_2 9.241569
Rin86_3 in86_2 in86_3 9.241569
Rin86_4 in86_3 in86_4 9.241569
Rin86_5 in86_4 in86_5 9.241569
Rin86_6 in86_5 in86_6 9.241569
Rin86_7 in86_6 in86_7 9.241569
Rin86_8 in86_7 in86_8 9.241569
Rin86_9 in86_8 in86_9 9.241569
Rin86_10 in86_9 in86_10 9.241569
Rin86_11 in86_10 in86_11 9.241569
Rin86_12 in86_11 in86_12 9.241569
Rin86_13 in86_12 in86_13 9.241569
Rin86_14 in86_13 in86_14 9.241569
Rin86_15 in86_14 in86_15 9.241569
Rin86_16 in86_15 in86_16 9.241569
Rin86_17 in86_16 in86_17 9.241569
Rin86_18 in86_17 in86_18 9.241569
Rin86_19 in86_18 in86_19 9.241569
Rin86_20 in86_19 in86_20 9.241569
Rin86_21 in86_20 in86_21 9.241569
Rin86_22 in86_21 in86_22 9.241569
Rin86_23 in86_22 in86_23 9.241569
Rin86_24 in86_23 in86_24 9.241569
Rin86_25 in86_24 in86_25 9.241569
Rin86_26 in86_25 in86_26 9.241569
Rin86_27 in86_26 in86_27 9.241569
Rin86_28 in86_27 in86_28 9.241569
Rin86_29 in86 in86_29 9.241569
Rin86_30 in86_29 in86_30 9.241569
Rin86_31 in86_30 in86_31 9.241569
Rin86_32 in86_31 in86_32 9.241569
Rin86_33 in86_32 in86_33 9.241569
Rin86_34 in86_33 in86_34 9.241569
Rin86_35 in86_34 in86_35 9.241569
Rin86_36 in86_35 in86_36 9.241569
Rin86_37 in86_36 in86_37 9.241569
Rin86_38 in86_37 in86_38 9.241569
Rin86_39 in86_38 in86_39 9.241569
Rin86_40 in86_39 in86_40 9.241569
Rin86_41 in86_40 in86_41 9.241569
Rin86_42 in86_41 in86_42 9.241569
Rin86_43 in86_42 in86_43 9.241569
Rin86_44 in86_43 in86_44 9.241569
Rin86_45 in86_44 in86_45 9.241569
Rin86_46 in86_45 in86_46 9.241569
Rin86_47 in86_46 in86_47 9.241569
Rin86_48 in86_47 in86_48 9.241569
Rin86_49 in86_48 in86_49 9.241569
Rin86_50 in86_49 in86_50 9.241569
Rin86_51 in86_50 in86_51 9.241569
Rin86_52 in86_51 in86_52 9.241569
Rin86_53 in86_52 in86_53 9.241569
Rin86_54 in86_53 in86_54 9.241569
Rin86_55 in86_54 in86_55 9.241569
Rin86_56 in86_55 in86_56 9.241569
Rin86_57 in86 in86_57 9.241569
Rin86_58 in86_57 in86_58 9.241569
Rin86_59 in86_58 in86_59 9.241569
Rin86_60 in86_59 in86_60 9.241569
Rin86_61 in86_60 in86_61 9.241569
Rin86_62 in86_61 in86_62 9.241569
Rin86_63 in86_62 in86_63 9.241569
Rin86_64 in86_63 in86_64 9.241569
Rin86_65 in86_64 in86_65 9.241569
Rin86_66 in86_65 in86_66 9.241569
Rin86_67 in86_66 in86_67 9.241569
Rin86_68 in86_67 in86_68 9.241569
Rin86_69 in86_68 in86_69 9.241569
Rin86_70 in86_69 in86_70 9.241569
Rin86_71 in86_70 in86_71 9.241569
Rin86_72 in86_71 in86_72 9.241569
Rin86_73 in86_72 in86_73 9.241569
Rin86_74 in86_73 in86_74 9.241569
Rin86_75 in86_74 in86_75 9.241569
Rin86_76 in86_75 in86_76 9.241569
Rin86_77 in86_76 in86_77 9.241569
Rin86_78 in86_77 in86_78 9.241569
Rin86_79 in86_78 in86_79 9.241569
Rin86_80 in86_79 in86_80 9.241569
Rin86_81 in86_80 in86_81 9.241569
Rin86_82 in86_81 in86_82 9.241569
Rin86_83 in86_82 in86_83 9.241569
Rin86_84 in86_83 in86_84 9.241569
Rin87_1 in87 in87_1 9.241569
Rin87_2 in87_1 in87_2 9.241569
Rin87_3 in87_2 in87_3 9.241569
Rin87_4 in87_3 in87_4 9.241569
Rin87_5 in87_4 in87_5 9.241569
Rin87_6 in87_5 in87_6 9.241569
Rin87_7 in87_6 in87_7 9.241569
Rin87_8 in87_7 in87_8 9.241569
Rin87_9 in87_8 in87_9 9.241569
Rin87_10 in87_9 in87_10 9.241569
Rin87_11 in87_10 in87_11 9.241569
Rin87_12 in87_11 in87_12 9.241569
Rin87_13 in87_12 in87_13 9.241569
Rin87_14 in87_13 in87_14 9.241569
Rin87_15 in87_14 in87_15 9.241569
Rin87_16 in87_15 in87_16 9.241569
Rin87_17 in87_16 in87_17 9.241569
Rin87_18 in87_17 in87_18 9.241569
Rin87_19 in87_18 in87_19 9.241569
Rin87_20 in87_19 in87_20 9.241569
Rin87_21 in87_20 in87_21 9.241569
Rin87_22 in87_21 in87_22 9.241569
Rin87_23 in87_22 in87_23 9.241569
Rin87_24 in87_23 in87_24 9.241569
Rin87_25 in87_24 in87_25 9.241569
Rin87_26 in87_25 in87_26 9.241569
Rin87_27 in87_26 in87_27 9.241569
Rin87_28 in87_27 in87_28 9.241569
Rin87_29 in87 in87_29 9.241569
Rin87_30 in87_29 in87_30 9.241569
Rin87_31 in87_30 in87_31 9.241569
Rin87_32 in87_31 in87_32 9.241569
Rin87_33 in87_32 in87_33 9.241569
Rin87_34 in87_33 in87_34 9.241569
Rin87_35 in87_34 in87_35 9.241569
Rin87_36 in87_35 in87_36 9.241569
Rin87_37 in87_36 in87_37 9.241569
Rin87_38 in87_37 in87_38 9.241569
Rin87_39 in87_38 in87_39 9.241569
Rin87_40 in87_39 in87_40 9.241569
Rin87_41 in87_40 in87_41 9.241569
Rin87_42 in87_41 in87_42 9.241569
Rin87_43 in87_42 in87_43 9.241569
Rin87_44 in87_43 in87_44 9.241569
Rin87_45 in87_44 in87_45 9.241569
Rin87_46 in87_45 in87_46 9.241569
Rin87_47 in87_46 in87_47 9.241569
Rin87_48 in87_47 in87_48 9.241569
Rin87_49 in87_48 in87_49 9.241569
Rin87_50 in87_49 in87_50 9.241569
Rin87_51 in87_50 in87_51 9.241569
Rin87_52 in87_51 in87_52 9.241569
Rin87_53 in87_52 in87_53 9.241569
Rin87_54 in87_53 in87_54 9.241569
Rin87_55 in87_54 in87_55 9.241569
Rin87_56 in87_55 in87_56 9.241569
Rin87_57 in87 in87_57 9.241569
Rin87_58 in87_57 in87_58 9.241569
Rin87_59 in87_58 in87_59 9.241569
Rin87_60 in87_59 in87_60 9.241569
Rin87_61 in87_60 in87_61 9.241569
Rin87_62 in87_61 in87_62 9.241569
Rin87_63 in87_62 in87_63 9.241569
Rin87_64 in87_63 in87_64 9.241569
Rin87_65 in87_64 in87_65 9.241569
Rin87_66 in87_65 in87_66 9.241569
Rin87_67 in87_66 in87_67 9.241569
Rin87_68 in87_67 in87_68 9.241569
Rin87_69 in87_68 in87_69 9.241569
Rin87_70 in87_69 in87_70 9.241569
Rin87_71 in87_70 in87_71 9.241569
Rin87_72 in87_71 in87_72 9.241569
Rin87_73 in87_72 in87_73 9.241569
Rin87_74 in87_73 in87_74 9.241569
Rin87_75 in87_74 in87_75 9.241569
Rin87_76 in87_75 in87_76 9.241569
Rin87_77 in87_76 in87_77 9.241569
Rin87_78 in87_77 in87_78 9.241569
Rin87_79 in87_78 in87_79 9.241569
Rin87_80 in87_79 in87_80 9.241569
Rin87_81 in87_80 in87_81 9.241569
Rin87_82 in87_81 in87_82 9.241569
Rin87_83 in87_82 in87_83 9.241569
Rin87_84 in87_83 in87_84 9.241569
Rin88_1 in88 in88_1 9.241569
Rin88_2 in88_1 in88_2 9.241569
Rin88_3 in88_2 in88_3 9.241569
Rin88_4 in88_3 in88_4 9.241569
Rin88_5 in88_4 in88_5 9.241569
Rin88_6 in88_5 in88_6 9.241569
Rin88_7 in88_6 in88_7 9.241569
Rin88_8 in88_7 in88_8 9.241569
Rin88_9 in88_8 in88_9 9.241569
Rin88_10 in88_9 in88_10 9.241569
Rin88_11 in88_10 in88_11 9.241569
Rin88_12 in88_11 in88_12 9.241569
Rin88_13 in88_12 in88_13 9.241569
Rin88_14 in88_13 in88_14 9.241569
Rin88_15 in88_14 in88_15 9.241569
Rin88_16 in88_15 in88_16 9.241569
Rin88_17 in88_16 in88_17 9.241569
Rin88_18 in88_17 in88_18 9.241569
Rin88_19 in88_18 in88_19 9.241569
Rin88_20 in88_19 in88_20 9.241569
Rin88_21 in88_20 in88_21 9.241569
Rin88_22 in88_21 in88_22 9.241569
Rin88_23 in88_22 in88_23 9.241569
Rin88_24 in88_23 in88_24 9.241569
Rin88_25 in88_24 in88_25 9.241569
Rin88_26 in88_25 in88_26 9.241569
Rin88_27 in88_26 in88_27 9.241569
Rin88_28 in88_27 in88_28 9.241569
Rin88_29 in88 in88_29 9.241569
Rin88_30 in88_29 in88_30 9.241569
Rin88_31 in88_30 in88_31 9.241569
Rin88_32 in88_31 in88_32 9.241569
Rin88_33 in88_32 in88_33 9.241569
Rin88_34 in88_33 in88_34 9.241569
Rin88_35 in88_34 in88_35 9.241569
Rin88_36 in88_35 in88_36 9.241569
Rin88_37 in88_36 in88_37 9.241569
Rin88_38 in88_37 in88_38 9.241569
Rin88_39 in88_38 in88_39 9.241569
Rin88_40 in88_39 in88_40 9.241569
Rin88_41 in88_40 in88_41 9.241569
Rin88_42 in88_41 in88_42 9.241569
Rin88_43 in88_42 in88_43 9.241569
Rin88_44 in88_43 in88_44 9.241569
Rin88_45 in88_44 in88_45 9.241569
Rin88_46 in88_45 in88_46 9.241569
Rin88_47 in88_46 in88_47 9.241569
Rin88_48 in88_47 in88_48 9.241569
Rin88_49 in88_48 in88_49 9.241569
Rin88_50 in88_49 in88_50 9.241569
Rin88_51 in88_50 in88_51 9.241569
Rin88_52 in88_51 in88_52 9.241569
Rin88_53 in88_52 in88_53 9.241569
Rin88_54 in88_53 in88_54 9.241569
Rin88_55 in88_54 in88_55 9.241569
Rin88_56 in88_55 in88_56 9.241569
Rin88_57 in88 in88_57 9.241569
Rin88_58 in88_57 in88_58 9.241569
Rin88_59 in88_58 in88_59 9.241569
Rin88_60 in88_59 in88_60 9.241569
Rin88_61 in88_60 in88_61 9.241569
Rin88_62 in88_61 in88_62 9.241569
Rin88_63 in88_62 in88_63 9.241569
Rin88_64 in88_63 in88_64 9.241569
Rin88_65 in88_64 in88_65 9.241569
Rin88_66 in88_65 in88_66 9.241569
Rin88_67 in88_66 in88_67 9.241569
Rin88_68 in88_67 in88_68 9.241569
Rin88_69 in88_68 in88_69 9.241569
Rin88_70 in88_69 in88_70 9.241569
Rin88_71 in88_70 in88_71 9.241569
Rin88_72 in88_71 in88_72 9.241569
Rin88_73 in88_72 in88_73 9.241569
Rin88_74 in88_73 in88_74 9.241569
Rin88_75 in88_74 in88_75 9.241569
Rin88_76 in88_75 in88_76 9.241569
Rin88_77 in88_76 in88_77 9.241569
Rin88_78 in88_77 in88_78 9.241569
Rin88_79 in88_78 in88_79 9.241569
Rin88_80 in88_79 in88_80 9.241569
Rin88_81 in88_80 in88_81 9.241569
Rin88_82 in88_81 in88_82 9.241569
Rin88_83 in88_82 in88_83 9.241569
Rin88_84 in88_83 in88_84 9.241569
Rin89_1 in89 in89_1 9.241569
Rin89_2 in89_1 in89_2 9.241569
Rin89_3 in89_2 in89_3 9.241569
Rin89_4 in89_3 in89_4 9.241569
Rin89_5 in89_4 in89_5 9.241569
Rin89_6 in89_5 in89_6 9.241569
Rin89_7 in89_6 in89_7 9.241569
Rin89_8 in89_7 in89_8 9.241569
Rin89_9 in89_8 in89_9 9.241569
Rin89_10 in89_9 in89_10 9.241569
Rin89_11 in89_10 in89_11 9.241569
Rin89_12 in89_11 in89_12 9.241569
Rin89_13 in89_12 in89_13 9.241569
Rin89_14 in89_13 in89_14 9.241569
Rin89_15 in89_14 in89_15 9.241569
Rin89_16 in89_15 in89_16 9.241569
Rin89_17 in89_16 in89_17 9.241569
Rin89_18 in89_17 in89_18 9.241569
Rin89_19 in89_18 in89_19 9.241569
Rin89_20 in89_19 in89_20 9.241569
Rin89_21 in89_20 in89_21 9.241569
Rin89_22 in89_21 in89_22 9.241569
Rin89_23 in89_22 in89_23 9.241569
Rin89_24 in89_23 in89_24 9.241569
Rin89_25 in89_24 in89_25 9.241569
Rin89_26 in89_25 in89_26 9.241569
Rin89_27 in89_26 in89_27 9.241569
Rin89_28 in89_27 in89_28 9.241569
Rin89_29 in89 in89_29 9.241569
Rin89_30 in89_29 in89_30 9.241569
Rin89_31 in89_30 in89_31 9.241569
Rin89_32 in89_31 in89_32 9.241569
Rin89_33 in89_32 in89_33 9.241569
Rin89_34 in89_33 in89_34 9.241569
Rin89_35 in89_34 in89_35 9.241569
Rin89_36 in89_35 in89_36 9.241569
Rin89_37 in89_36 in89_37 9.241569
Rin89_38 in89_37 in89_38 9.241569
Rin89_39 in89_38 in89_39 9.241569
Rin89_40 in89_39 in89_40 9.241569
Rin89_41 in89_40 in89_41 9.241569
Rin89_42 in89_41 in89_42 9.241569
Rin89_43 in89_42 in89_43 9.241569
Rin89_44 in89_43 in89_44 9.241569
Rin89_45 in89_44 in89_45 9.241569
Rin89_46 in89_45 in89_46 9.241569
Rin89_47 in89_46 in89_47 9.241569
Rin89_48 in89_47 in89_48 9.241569
Rin89_49 in89_48 in89_49 9.241569
Rin89_50 in89_49 in89_50 9.241569
Rin89_51 in89_50 in89_51 9.241569
Rin89_52 in89_51 in89_52 9.241569
Rin89_53 in89_52 in89_53 9.241569
Rin89_54 in89_53 in89_54 9.241569
Rin89_55 in89_54 in89_55 9.241569
Rin89_56 in89_55 in89_56 9.241569
Rin89_57 in89 in89_57 9.241569
Rin89_58 in89_57 in89_58 9.241569
Rin89_59 in89_58 in89_59 9.241569
Rin89_60 in89_59 in89_60 9.241569
Rin89_61 in89_60 in89_61 9.241569
Rin89_62 in89_61 in89_62 9.241569
Rin89_63 in89_62 in89_63 9.241569
Rin89_64 in89_63 in89_64 9.241569
Rin89_65 in89_64 in89_65 9.241569
Rin89_66 in89_65 in89_66 9.241569
Rin89_67 in89_66 in89_67 9.241569
Rin89_68 in89_67 in89_68 9.241569
Rin89_69 in89_68 in89_69 9.241569
Rin89_70 in89_69 in89_70 9.241569
Rin89_71 in89_70 in89_71 9.241569
Rin89_72 in89_71 in89_72 9.241569
Rin89_73 in89_72 in89_73 9.241569
Rin89_74 in89_73 in89_74 9.241569
Rin89_75 in89_74 in89_75 9.241569
Rin89_76 in89_75 in89_76 9.241569
Rin89_77 in89_76 in89_77 9.241569
Rin89_78 in89_77 in89_78 9.241569
Rin89_79 in89_78 in89_79 9.241569
Rin89_80 in89_79 in89_80 9.241569
Rin89_81 in89_80 in89_81 9.241569
Rin89_82 in89_81 in89_82 9.241569
Rin89_83 in89_82 in89_83 9.241569
Rin89_84 in89_83 in89_84 9.241569
Rin90_1 in90 in90_1 9.241569
Rin90_2 in90_1 in90_2 9.241569
Rin90_3 in90_2 in90_3 9.241569
Rin90_4 in90_3 in90_4 9.241569
Rin90_5 in90_4 in90_5 9.241569
Rin90_6 in90_5 in90_6 9.241569
Rin90_7 in90_6 in90_7 9.241569
Rin90_8 in90_7 in90_8 9.241569
Rin90_9 in90_8 in90_9 9.241569
Rin90_10 in90_9 in90_10 9.241569
Rin90_11 in90_10 in90_11 9.241569
Rin90_12 in90_11 in90_12 9.241569
Rin90_13 in90_12 in90_13 9.241569
Rin90_14 in90_13 in90_14 9.241569
Rin90_15 in90_14 in90_15 9.241569
Rin90_16 in90_15 in90_16 9.241569
Rin90_17 in90_16 in90_17 9.241569
Rin90_18 in90_17 in90_18 9.241569
Rin90_19 in90_18 in90_19 9.241569
Rin90_20 in90_19 in90_20 9.241569
Rin90_21 in90_20 in90_21 9.241569
Rin90_22 in90_21 in90_22 9.241569
Rin90_23 in90_22 in90_23 9.241569
Rin90_24 in90_23 in90_24 9.241569
Rin90_25 in90_24 in90_25 9.241569
Rin90_26 in90_25 in90_26 9.241569
Rin90_27 in90_26 in90_27 9.241569
Rin90_28 in90_27 in90_28 9.241569
Rin90_29 in90 in90_29 9.241569
Rin90_30 in90_29 in90_30 9.241569
Rin90_31 in90_30 in90_31 9.241569
Rin90_32 in90_31 in90_32 9.241569
Rin90_33 in90_32 in90_33 9.241569
Rin90_34 in90_33 in90_34 9.241569
Rin90_35 in90_34 in90_35 9.241569
Rin90_36 in90_35 in90_36 9.241569
Rin90_37 in90_36 in90_37 9.241569
Rin90_38 in90_37 in90_38 9.241569
Rin90_39 in90_38 in90_39 9.241569
Rin90_40 in90_39 in90_40 9.241569
Rin90_41 in90_40 in90_41 9.241569
Rin90_42 in90_41 in90_42 9.241569
Rin90_43 in90_42 in90_43 9.241569
Rin90_44 in90_43 in90_44 9.241569
Rin90_45 in90_44 in90_45 9.241569
Rin90_46 in90_45 in90_46 9.241569
Rin90_47 in90_46 in90_47 9.241569
Rin90_48 in90_47 in90_48 9.241569
Rin90_49 in90_48 in90_49 9.241569
Rin90_50 in90_49 in90_50 9.241569
Rin90_51 in90_50 in90_51 9.241569
Rin90_52 in90_51 in90_52 9.241569
Rin90_53 in90_52 in90_53 9.241569
Rin90_54 in90_53 in90_54 9.241569
Rin90_55 in90_54 in90_55 9.241569
Rin90_56 in90_55 in90_56 9.241569
Rin90_57 in90 in90_57 9.241569
Rin90_58 in90_57 in90_58 9.241569
Rin90_59 in90_58 in90_59 9.241569
Rin90_60 in90_59 in90_60 9.241569
Rin90_61 in90_60 in90_61 9.241569
Rin90_62 in90_61 in90_62 9.241569
Rin90_63 in90_62 in90_63 9.241569
Rin90_64 in90_63 in90_64 9.241569
Rin90_65 in90_64 in90_65 9.241569
Rin90_66 in90_65 in90_66 9.241569
Rin90_67 in90_66 in90_67 9.241569
Rin90_68 in90_67 in90_68 9.241569
Rin90_69 in90_68 in90_69 9.241569
Rin90_70 in90_69 in90_70 9.241569
Rin90_71 in90_70 in90_71 9.241569
Rin90_72 in90_71 in90_72 9.241569
Rin90_73 in90_72 in90_73 9.241569
Rin90_74 in90_73 in90_74 9.241569
Rin90_75 in90_74 in90_75 9.241569
Rin90_76 in90_75 in90_76 9.241569
Rin90_77 in90_76 in90_77 9.241569
Rin90_78 in90_77 in90_78 9.241569
Rin90_79 in90_78 in90_79 9.241569
Rin90_80 in90_79 in90_80 9.241569
Rin90_81 in90_80 in90_81 9.241569
Rin90_82 in90_81 in90_82 9.241569
Rin90_83 in90_82 in90_83 9.241569
Rin90_84 in90_83 in90_84 9.241569
Rin91_1 in91 in91_1 9.241569
Rin91_2 in91_1 in91_2 9.241569
Rin91_3 in91_2 in91_3 9.241569
Rin91_4 in91_3 in91_4 9.241569
Rin91_5 in91_4 in91_5 9.241569
Rin91_6 in91_5 in91_6 9.241569
Rin91_7 in91_6 in91_7 9.241569
Rin91_8 in91_7 in91_8 9.241569
Rin91_9 in91_8 in91_9 9.241569
Rin91_10 in91_9 in91_10 9.241569
Rin91_11 in91_10 in91_11 9.241569
Rin91_12 in91_11 in91_12 9.241569
Rin91_13 in91_12 in91_13 9.241569
Rin91_14 in91_13 in91_14 9.241569
Rin91_15 in91_14 in91_15 9.241569
Rin91_16 in91_15 in91_16 9.241569
Rin91_17 in91_16 in91_17 9.241569
Rin91_18 in91_17 in91_18 9.241569
Rin91_19 in91_18 in91_19 9.241569
Rin91_20 in91_19 in91_20 9.241569
Rin91_21 in91_20 in91_21 9.241569
Rin91_22 in91_21 in91_22 9.241569
Rin91_23 in91_22 in91_23 9.241569
Rin91_24 in91_23 in91_24 9.241569
Rin91_25 in91_24 in91_25 9.241569
Rin91_26 in91_25 in91_26 9.241569
Rin91_27 in91_26 in91_27 9.241569
Rin91_28 in91_27 in91_28 9.241569
Rin91_29 in91 in91_29 9.241569
Rin91_30 in91_29 in91_30 9.241569
Rin91_31 in91_30 in91_31 9.241569
Rin91_32 in91_31 in91_32 9.241569
Rin91_33 in91_32 in91_33 9.241569
Rin91_34 in91_33 in91_34 9.241569
Rin91_35 in91_34 in91_35 9.241569
Rin91_36 in91_35 in91_36 9.241569
Rin91_37 in91_36 in91_37 9.241569
Rin91_38 in91_37 in91_38 9.241569
Rin91_39 in91_38 in91_39 9.241569
Rin91_40 in91_39 in91_40 9.241569
Rin91_41 in91_40 in91_41 9.241569
Rin91_42 in91_41 in91_42 9.241569
Rin91_43 in91_42 in91_43 9.241569
Rin91_44 in91_43 in91_44 9.241569
Rin91_45 in91_44 in91_45 9.241569
Rin91_46 in91_45 in91_46 9.241569
Rin91_47 in91_46 in91_47 9.241569
Rin91_48 in91_47 in91_48 9.241569
Rin91_49 in91_48 in91_49 9.241569
Rin91_50 in91_49 in91_50 9.241569
Rin91_51 in91_50 in91_51 9.241569
Rin91_52 in91_51 in91_52 9.241569
Rin91_53 in91_52 in91_53 9.241569
Rin91_54 in91_53 in91_54 9.241569
Rin91_55 in91_54 in91_55 9.241569
Rin91_56 in91_55 in91_56 9.241569
Rin91_57 in91 in91_57 9.241569
Rin91_58 in91_57 in91_58 9.241569
Rin91_59 in91_58 in91_59 9.241569
Rin91_60 in91_59 in91_60 9.241569
Rin91_61 in91_60 in91_61 9.241569
Rin91_62 in91_61 in91_62 9.241569
Rin91_63 in91_62 in91_63 9.241569
Rin91_64 in91_63 in91_64 9.241569
Rin91_65 in91_64 in91_65 9.241569
Rin91_66 in91_65 in91_66 9.241569
Rin91_67 in91_66 in91_67 9.241569
Rin91_68 in91_67 in91_68 9.241569
Rin91_69 in91_68 in91_69 9.241569
Rin91_70 in91_69 in91_70 9.241569
Rin91_71 in91_70 in91_71 9.241569
Rin91_72 in91_71 in91_72 9.241569
Rin91_73 in91_72 in91_73 9.241569
Rin91_74 in91_73 in91_74 9.241569
Rin91_75 in91_74 in91_75 9.241569
Rin91_76 in91_75 in91_76 9.241569
Rin91_77 in91_76 in91_77 9.241569
Rin91_78 in91_77 in91_78 9.241569
Rin91_79 in91_78 in91_79 9.241569
Rin91_80 in91_79 in91_80 9.241569
Rin91_81 in91_80 in91_81 9.241569
Rin91_82 in91_81 in91_82 9.241569
Rin91_83 in91_82 in91_83 9.241569
Rin91_84 in91_83 in91_84 9.241569
Rin92_1 in92 in92_1 9.241569
Rin92_2 in92_1 in92_2 9.241569
Rin92_3 in92_2 in92_3 9.241569
Rin92_4 in92_3 in92_4 9.241569
Rin92_5 in92_4 in92_5 9.241569
Rin92_6 in92_5 in92_6 9.241569
Rin92_7 in92_6 in92_7 9.241569
Rin92_8 in92_7 in92_8 9.241569
Rin92_9 in92_8 in92_9 9.241569
Rin92_10 in92_9 in92_10 9.241569
Rin92_11 in92_10 in92_11 9.241569
Rin92_12 in92_11 in92_12 9.241569
Rin92_13 in92_12 in92_13 9.241569
Rin92_14 in92_13 in92_14 9.241569
Rin92_15 in92_14 in92_15 9.241569
Rin92_16 in92_15 in92_16 9.241569
Rin92_17 in92_16 in92_17 9.241569
Rin92_18 in92_17 in92_18 9.241569
Rin92_19 in92_18 in92_19 9.241569
Rin92_20 in92_19 in92_20 9.241569
Rin92_21 in92_20 in92_21 9.241569
Rin92_22 in92_21 in92_22 9.241569
Rin92_23 in92_22 in92_23 9.241569
Rin92_24 in92_23 in92_24 9.241569
Rin92_25 in92_24 in92_25 9.241569
Rin92_26 in92_25 in92_26 9.241569
Rin92_27 in92_26 in92_27 9.241569
Rin92_28 in92_27 in92_28 9.241569
Rin92_29 in92 in92_29 9.241569
Rin92_30 in92_29 in92_30 9.241569
Rin92_31 in92_30 in92_31 9.241569
Rin92_32 in92_31 in92_32 9.241569
Rin92_33 in92_32 in92_33 9.241569
Rin92_34 in92_33 in92_34 9.241569
Rin92_35 in92_34 in92_35 9.241569
Rin92_36 in92_35 in92_36 9.241569
Rin92_37 in92_36 in92_37 9.241569
Rin92_38 in92_37 in92_38 9.241569
Rin92_39 in92_38 in92_39 9.241569
Rin92_40 in92_39 in92_40 9.241569
Rin92_41 in92_40 in92_41 9.241569
Rin92_42 in92_41 in92_42 9.241569
Rin92_43 in92_42 in92_43 9.241569
Rin92_44 in92_43 in92_44 9.241569
Rin92_45 in92_44 in92_45 9.241569
Rin92_46 in92_45 in92_46 9.241569
Rin92_47 in92_46 in92_47 9.241569
Rin92_48 in92_47 in92_48 9.241569
Rin92_49 in92_48 in92_49 9.241569
Rin92_50 in92_49 in92_50 9.241569
Rin92_51 in92_50 in92_51 9.241569
Rin92_52 in92_51 in92_52 9.241569
Rin92_53 in92_52 in92_53 9.241569
Rin92_54 in92_53 in92_54 9.241569
Rin92_55 in92_54 in92_55 9.241569
Rin92_56 in92_55 in92_56 9.241569
Rin92_57 in92 in92_57 9.241569
Rin92_58 in92_57 in92_58 9.241569
Rin92_59 in92_58 in92_59 9.241569
Rin92_60 in92_59 in92_60 9.241569
Rin92_61 in92_60 in92_61 9.241569
Rin92_62 in92_61 in92_62 9.241569
Rin92_63 in92_62 in92_63 9.241569
Rin92_64 in92_63 in92_64 9.241569
Rin92_65 in92_64 in92_65 9.241569
Rin92_66 in92_65 in92_66 9.241569
Rin92_67 in92_66 in92_67 9.241569
Rin92_68 in92_67 in92_68 9.241569
Rin92_69 in92_68 in92_69 9.241569
Rin92_70 in92_69 in92_70 9.241569
Rin92_71 in92_70 in92_71 9.241569
Rin92_72 in92_71 in92_72 9.241569
Rin92_73 in92_72 in92_73 9.241569
Rin92_74 in92_73 in92_74 9.241569
Rin92_75 in92_74 in92_75 9.241569
Rin92_76 in92_75 in92_76 9.241569
Rin92_77 in92_76 in92_77 9.241569
Rin92_78 in92_77 in92_78 9.241569
Rin92_79 in92_78 in92_79 9.241569
Rin92_80 in92_79 in92_80 9.241569
Rin92_81 in92_80 in92_81 9.241569
Rin92_82 in92_81 in92_82 9.241569
Rin92_83 in92_82 in92_83 9.241569
Rin92_84 in92_83 in92_84 9.241569
Rin93_1 in93 in93_1 9.241569
Rin93_2 in93_1 in93_2 9.241569
Rin93_3 in93_2 in93_3 9.241569
Rin93_4 in93_3 in93_4 9.241569
Rin93_5 in93_4 in93_5 9.241569
Rin93_6 in93_5 in93_6 9.241569
Rin93_7 in93_6 in93_7 9.241569
Rin93_8 in93_7 in93_8 9.241569
Rin93_9 in93_8 in93_9 9.241569
Rin93_10 in93_9 in93_10 9.241569
Rin93_11 in93_10 in93_11 9.241569
Rin93_12 in93_11 in93_12 9.241569
Rin93_13 in93_12 in93_13 9.241569
Rin93_14 in93_13 in93_14 9.241569
Rin93_15 in93_14 in93_15 9.241569
Rin93_16 in93_15 in93_16 9.241569
Rin93_17 in93_16 in93_17 9.241569
Rin93_18 in93_17 in93_18 9.241569
Rin93_19 in93_18 in93_19 9.241569
Rin93_20 in93_19 in93_20 9.241569
Rin93_21 in93_20 in93_21 9.241569
Rin93_22 in93_21 in93_22 9.241569
Rin93_23 in93_22 in93_23 9.241569
Rin93_24 in93_23 in93_24 9.241569
Rin93_25 in93_24 in93_25 9.241569
Rin93_26 in93_25 in93_26 9.241569
Rin93_27 in93_26 in93_27 9.241569
Rin93_28 in93_27 in93_28 9.241569
Rin93_29 in93 in93_29 9.241569
Rin93_30 in93_29 in93_30 9.241569
Rin93_31 in93_30 in93_31 9.241569
Rin93_32 in93_31 in93_32 9.241569
Rin93_33 in93_32 in93_33 9.241569
Rin93_34 in93_33 in93_34 9.241569
Rin93_35 in93_34 in93_35 9.241569
Rin93_36 in93_35 in93_36 9.241569
Rin93_37 in93_36 in93_37 9.241569
Rin93_38 in93_37 in93_38 9.241569
Rin93_39 in93_38 in93_39 9.241569
Rin93_40 in93_39 in93_40 9.241569
Rin93_41 in93_40 in93_41 9.241569
Rin93_42 in93_41 in93_42 9.241569
Rin93_43 in93_42 in93_43 9.241569
Rin93_44 in93_43 in93_44 9.241569
Rin93_45 in93_44 in93_45 9.241569
Rin93_46 in93_45 in93_46 9.241569
Rin93_47 in93_46 in93_47 9.241569
Rin93_48 in93_47 in93_48 9.241569
Rin93_49 in93_48 in93_49 9.241569
Rin93_50 in93_49 in93_50 9.241569
Rin93_51 in93_50 in93_51 9.241569
Rin93_52 in93_51 in93_52 9.241569
Rin93_53 in93_52 in93_53 9.241569
Rin93_54 in93_53 in93_54 9.241569
Rin93_55 in93_54 in93_55 9.241569
Rin93_56 in93_55 in93_56 9.241569
Rin93_57 in93 in93_57 9.241569
Rin93_58 in93_57 in93_58 9.241569
Rin93_59 in93_58 in93_59 9.241569
Rin93_60 in93_59 in93_60 9.241569
Rin93_61 in93_60 in93_61 9.241569
Rin93_62 in93_61 in93_62 9.241569
Rin93_63 in93_62 in93_63 9.241569
Rin93_64 in93_63 in93_64 9.241569
Rin93_65 in93_64 in93_65 9.241569
Rin93_66 in93_65 in93_66 9.241569
Rin93_67 in93_66 in93_67 9.241569
Rin93_68 in93_67 in93_68 9.241569
Rin93_69 in93_68 in93_69 9.241569
Rin93_70 in93_69 in93_70 9.241569
Rin93_71 in93_70 in93_71 9.241569
Rin93_72 in93_71 in93_72 9.241569
Rin93_73 in93_72 in93_73 9.241569
Rin93_74 in93_73 in93_74 9.241569
Rin93_75 in93_74 in93_75 9.241569
Rin93_76 in93_75 in93_76 9.241569
Rin93_77 in93_76 in93_77 9.241569
Rin93_78 in93_77 in93_78 9.241569
Rin93_79 in93_78 in93_79 9.241569
Rin93_80 in93_79 in93_80 9.241569
Rin93_81 in93_80 in93_81 9.241569
Rin93_82 in93_81 in93_82 9.241569
Rin93_83 in93_82 in93_83 9.241569
Rin93_84 in93_83 in93_84 9.241569
Rin94_1 in94 in94_1 9.241569
Rin94_2 in94_1 in94_2 9.241569
Rin94_3 in94_2 in94_3 9.241569
Rin94_4 in94_3 in94_4 9.241569
Rin94_5 in94_4 in94_5 9.241569
Rin94_6 in94_5 in94_6 9.241569
Rin94_7 in94_6 in94_7 9.241569
Rin94_8 in94_7 in94_8 9.241569
Rin94_9 in94_8 in94_9 9.241569
Rin94_10 in94_9 in94_10 9.241569
Rin94_11 in94_10 in94_11 9.241569
Rin94_12 in94_11 in94_12 9.241569
Rin94_13 in94_12 in94_13 9.241569
Rin94_14 in94_13 in94_14 9.241569
Rin94_15 in94_14 in94_15 9.241569
Rin94_16 in94_15 in94_16 9.241569
Rin94_17 in94_16 in94_17 9.241569
Rin94_18 in94_17 in94_18 9.241569
Rin94_19 in94_18 in94_19 9.241569
Rin94_20 in94_19 in94_20 9.241569
Rin94_21 in94_20 in94_21 9.241569
Rin94_22 in94_21 in94_22 9.241569
Rin94_23 in94_22 in94_23 9.241569
Rin94_24 in94_23 in94_24 9.241569
Rin94_25 in94_24 in94_25 9.241569
Rin94_26 in94_25 in94_26 9.241569
Rin94_27 in94_26 in94_27 9.241569
Rin94_28 in94_27 in94_28 9.241569
Rin94_29 in94 in94_29 9.241569
Rin94_30 in94_29 in94_30 9.241569
Rin94_31 in94_30 in94_31 9.241569
Rin94_32 in94_31 in94_32 9.241569
Rin94_33 in94_32 in94_33 9.241569
Rin94_34 in94_33 in94_34 9.241569
Rin94_35 in94_34 in94_35 9.241569
Rin94_36 in94_35 in94_36 9.241569
Rin94_37 in94_36 in94_37 9.241569
Rin94_38 in94_37 in94_38 9.241569
Rin94_39 in94_38 in94_39 9.241569
Rin94_40 in94_39 in94_40 9.241569
Rin94_41 in94_40 in94_41 9.241569
Rin94_42 in94_41 in94_42 9.241569
Rin94_43 in94_42 in94_43 9.241569
Rin94_44 in94_43 in94_44 9.241569
Rin94_45 in94_44 in94_45 9.241569
Rin94_46 in94_45 in94_46 9.241569
Rin94_47 in94_46 in94_47 9.241569
Rin94_48 in94_47 in94_48 9.241569
Rin94_49 in94_48 in94_49 9.241569
Rin94_50 in94_49 in94_50 9.241569
Rin94_51 in94_50 in94_51 9.241569
Rin94_52 in94_51 in94_52 9.241569
Rin94_53 in94_52 in94_53 9.241569
Rin94_54 in94_53 in94_54 9.241569
Rin94_55 in94_54 in94_55 9.241569
Rin94_56 in94_55 in94_56 9.241569
Rin94_57 in94 in94_57 9.241569
Rin94_58 in94_57 in94_58 9.241569
Rin94_59 in94_58 in94_59 9.241569
Rin94_60 in94_59 in94_60 9.241569
Rin94_61 in94_60 in94_61 9.241569
Rin94_62 in94_61 in94_62 9.241569
Rin94_63 in94_62 in94_63 9.241569
Rin94_64 in94_63 in94_64 9.241569
Rin94_65 in94_64 in94_65 9.241569
Rin94_66 in94_65 in94_66 9.241569
Rin94_67 in94_66 in94_67 9.241569
Rin94_68 in94_67 in94_68 9.241569
Rin94_69 in94_68 in94_69 9.241569
Rin94_70 in94_69 in94_70 9.241569
Rin94_71 in94_70 in94_71 9.241569
Rin94_72 in94_71 in94_72 9.241569
Rin94_73 in94_72 in94_73 9.241569
Rin94_74 in94_73 in94_74 9.241569
Rin94_75 in94_74 in94_75 9.241569
Rin94_76 in94_75 in94_76 9.241569
Rin94_77 in94_76 in94_77 9.241569
Rin94_78 in94_77 in94_78 9.241569
Rin94_79 in94_78 in94_79 9.241569
Rin94_80 in94_79 in94_80 9.241569
Rin94_81 in94_80 in94_81 9.241569
Rin94_82 in94_81 in94_82 9.241569
Rin94_83 in94_82 in94_83 9.241569
Rin94_84 in94_83 in94_84 9.241569
Rin95_1 in95 in95_1 9.241569
Rin95_2 in95_1 in95_2 9.241569
Rin95_3 in95_2 in95_3 9.241569
Rin95_4 in95_3 in95_4 9.241569
Rin95_5 in95_4 in95_5 9.241569
Rin95_6 in95_5 in95_6 9.241569
Rin95_7 in95_6 in95_7 9.241569
Rin95_8 in95_7 in95_8 9.241569
Rin95_9 in95_8 in95_9 9.241569
Rin95_10 in95_9 in95_10 9.241569
Rin95_11 in95_10 in95_11 9.241569
Rin95_12 in95_11 in95_12 9.241569
Rin95_13 in95_12 in95_13 9.241569
Rin95_14 in95_13 in95_14 9.241569
Rin95_15 in95_14 in95_15 9.241569
Rin95_16 in95_15 in95_16 9.241569
Rin95_17 in95_16 in95_17 9.241569
Rin95_18 in95_17 in95_18 9.241569
Rin95_19 in95_18 in95_19 9.241569
Rin95_20 in95_19 in95_20 9.241569
Rin95_21 in95_20 in95_21 9.241569
Rin95_22 in95_21 in95_22 9.241569
Rin95_23 in95_22 in95_23 9.241569
Rin95_24 in95_23 in95_24 9.241569
Rin95_25 in95_24 in95_25 9.241569
Rin95_26 in95_25 in95_26 9.241569
Rin95_27 in95_26 in95_27 9.241569
Rin95_28 in95_27 in95_28 9.241569
Rin95_29 in95 in95_29 9.241569
Rin95_30 in95_29 in95_30 9.241569
Rin95_31 in95_30 in95_31 9.241569
Rin95_32 in95_31 in95_32 9.241569
Rin95_33 in95_32 in95_33 9.241569
Rin95_34 in95_33 in95_34 9.241569
Rin95_35 in95_34 in95_35 9.241569
Rin95_36 in95_35 in95_36 9.241569
Rin95_37 in95_36 in95_37 9.241569
Rin95_38 in95_37 in95_38 9.241569
Rin95_39 in95_38 in95_39 9.241569
Rin95_40 in95_39 in95_40 9.241569
Rin95_41 in95_40 in95_41 9.241569
Rin95_42 in95_41 in95_42 9.241569
Rin95_43 in95_42 in95_43 9.241569
Rin95_44 in95_43 in95_44 9.241569
Rin95_45 in95_44 in95_45 9.241569
Rin95_46 in95_45 in95_46 9.241569
Rin95_47 in95_46 in95_47 9.241569
Rin95_48 in95_47 in95_48 9.241569
Rin95_49 in95_48 in95_49 9.241569
Rin95_50 in95_49 in95_50 9.241569
Rin95_51 in95_50 in95_51 9.241569
Rin95_52 in95_51 in95_52 9.241569
Rin95_53 in95_52 in95_53 9.241569
Rin95_54 in95_53 in95_54 9.241569
Rin95_55 in95_54 in95_55 9.241569
Rin95_56 in95_55 in95_56 9.241569
Rin95_57 in95 in95_57 9.241569
Rin95_58 in95_57 in95_58 9.241569
Rin95_59 in95_58 in95_59 9.241569
Rin95_60 in95_59 in95_60 9.241569
Rin95_61 in95_60 in95_61 9.241569
Rin95_62 in95_61 in95_62 9.241569
Rin95_63 in95_62 in95_63 9.241569
Rin95_64 in95_63 in95_64 9.241569
Rin95_65 in95_64 in95_65 9.241569
Rin95_66 in95_65 in95_66 9.241569
Rin95_67 in95_66 in95_67 9.241569
Rin95_68 in95_67 in95_68 9.241569
Rin95_69 in95_68 in95_69 9.241569
Rin95_70 in95_69 in95_70 9.241569
Rin95_71 in95_70 in95_71 9.241569
Rin95_72 in95_71 in95_72 9.241569
Rin95_73 in95_72 in95_73 9.241569
Rin95_74 in95_73 in95_74 9.241569
Rin95_75 in95_74 in95_75 9.241569
Rin95_76 in95_75 in95_76 9.241569
Rin95_77 in95_76 in95_77 9.241569
Rin95_78 in95_77 in95_78 9.241569
Rin95_79 in95_78 in95_79 9.241569
Rin95_80 in95_79 in95_80 9.241569
Rin95_81 in95_80 in95_81 9.241569
Rin95_82 in95_81 in95_82 9.241569
Rin95_83 in95_82 in95_83 9.241569
Rin95_84 in95_83 in95_84 9.241569
Rin96_1 in96 in96_1 9.241569
Rin96_2 in96_1 in96_2 9.241569
Rin96_3 in96_2 in96_3 9.241569
Rin96_4 in96_3 in96_4 9.241569
Rin96_5 in96_4 in96_5 9.241569
Rin96_6 in96_5 in96_6 9.241569
Rin96_7 in96_6 in96_7 9.241569
Rin96_8 in96_7 in96_8 9.241569
Rin96_9 in96_8 in96_9 9.241569
Rin96_10 in96_9 in96_10 9.241569
Rin96_11 in96_10 in96_11 9.241569
Rin96_12 in96_11 in96_12 9.241569
Rin96_13 in96_12 in96_13 9.241569
Rin96_14 in96_13 in96_14 9.241569
Rin96_15 in96_14 in96_15 9.241569
Rin96_16 in96_15 in96_16 9.241569
Rin96_17 in96_16 in96_17 9.241569
Rin96_18 in96_17 in96_18 9.241569
Rin96_19 in96_18 in96_19 9.241569
Rin96_20 in96_19 in96_20 9.241569
Rin96_21 in96_20 in96_21 9.241569
Rin96_22 in96_21 in96_22 9.241569
Rin96_23 in96_22 in96_23 9.241569
Rin96_24 in96_23 in96_24 9.241569
Rin96_25 in96_24 in96_25 9.241569
Rin96_26 in96_25 in96_26 9.241569
Rin96_27 in96_26 in96_27 9.241569
Rin96_28 in96_27 in96_28 9.241569
Rin96_29 in96 in96_29 9.241569
Rin96_30 in96_29 in96_30 9.241569
Rin96_31 in96_30 in96_31 9.241569
Rin96_32 in96_31 in96_32 9.241569
Rin96_33 in96_32 in96_33 9.241569
Rin96_34 in96_33 in96_34 9.241569
Rin96_35 in96_34 in96_35 9.241569
Rin96_36 in96_35 in96_36 9.241569
Rin96_37 in96_36 in96_37 9.241569
Rin96_38 in96_37 in96_38 9.241569
Rin96_39 in96_38 in96_39 9.241569
Rin96_40 in96_39 in96_40 9.241569
Rin96_41 in96_40 in96_41 9.241569
Rin96_42 in96_41 in96_42 9.241569
Rin96_43 in96_42 in96_43 9.241569
Rin96_44 in96_43 in96_44 9.241569
Rin96_45 in96_44 in96_45 9.241569
Rin96_46 in96_45 in96_46 9.241569
Rin96_47 in96_46 in96_47 9.241569
Rin96_48 in96_47 in96_48 9.241569
Rin96_49 in96_48 in96_49 9.241569
Rin96_50 in96_49 in96_50 9.241569
Rin96_51 in96_50 in96_51 9.241569
Rin96_52 in96_51 in96_52 9.241569
Rin96_53 in96_52 in96_53 9.241569
Rin96_54 in96_53 in96_54 9.241569
Rin96_55 in96_54 in96_55 9.241569
Rin96_56 in96_55 in96_56 9.241569
Rin96_57 in96 in96_57 9.241569
Rin96_58 in96_57 in96_58 9.241569
Rin96_59 in96_58 in96_59 9.241569
Rin96_60 in96_59 in96_60 9.241569
Rin96_61 in96_60 in96_61 9.241569
Rin96_62 in96_61 in96_62 9.241569
Rin96_63 in96_62 in96_63 9.241569
Rin96_64 in96_63 in96_64 9.241569
Rin96_65 in96_64 in96_65 9.241569
Rin96_66 in96_65 in96_66 9.241569
Rin96_67 in96_66 in96_67 9.241569
Rin96_68 in96_67 in96_68 9.241569
Rin96_69 in96_68 in96_69 9.241569
Rin96_70 in96_69 in96_70 9.241569
Rin96_71 in96_70 in96_71 9.241569
Rin96_72 in96_71 in96_72 9.241569
Rin96_73 in96_72 in96_73 9.241569
Rin96_74 in96_73 in96_74 9.241569
Rin96_75 in96_74 in96_75 9.241569
Rin96_76 in96_75 in96_76 9.241569
Rin96_77 in96_76 in96_77 9.241569
Rin96_78 in96_77 in96_78 9.241569
Rin96_79 in96_78 in96_79 9.241569
Rin96_80 in96_79 in96_80 9.241569
Rin96_81 in96_80 in96_81 9.241569
Rin96_82 in96_81 in96_82 9.241569
Rin96_83 in96_82 in96_83 9.241569
Rin96_84 in96_83 in96_84 9.241569
Rin97_1 in97 in97_1 9.241569
Rin97_2 in97_1 in97_2 9.241569
Rin97_3 in97_2 in97_3 9.241569
Rin97_4 in97_3 in97_4 9.241569
Rin97_5 in97_4 in97_5 9.241569
Rin97_6 in97_5 in97_6 9.241569
Rin97_7 in97_6 in97_7 9.241569
Rin97_8 in97_7 in97_8 9.241569
Rin97_9 in97_8 in97_9 9.241569
Rin97_10 in97_9 in97_10 9.241569
Rin97_11 in97_10 in97_11 9.241569
Rin97_12 in97_11 in97_12 9.241569
Rin97_13 in97_12 in97_13 9.241569
Rin97_14 in97_13 in97_14 9.241569
Rin97_15 in97_14 in97_15 9.241569
Rin97_16 in97_15 in97_16 9.241569
Rin97_17 in97_16 in97_17 9.241569
Rin97_18 in97_17 in97_18 9.241569
Rin97_19 in97_18 in97_19 9.241569
Rin97_20 in97_19 in97_20 9.241569
Rin97_21 in97_20 in97_21 9.241569
Rin97_22 in97_21 in97_22 9.241569
Rin97_23 in97_22 in97_23 9.241569
Rin97_24 in97_23 in97_24 9.241569
Rin97_25 in97_24 in97_25 9.241569
Rin97_26 in97_25 in97_26 9.241569
Rin97_27 in97_26 in97_27 9.241569
Rin97_28 in97_27 in97_28 9.241569
Rin97_29 in97 in97_29 9.241569
Rin97_30 in97_29 in97_30 9.241569
Rin97_31 in97_30 in97_31 9.241569
Rin97_32 in97_31 in97_32 9.241569
Rin97_33 in97_32 in97_33 9.241569
Rin97_34 in97_33 in97_34 9.241569
Rin97_35 in97_34 in97_35 9.241569
Rin97_36 in97_35 in97_36 9.241569
Rin97_37 in97_36 in97_37 9.241569
Rin97_38 in97_37 in97_38 9.241569
Rin97_39 in97_38 in97_39 9.241569
Rin97_40 in97_39 in97_40 9.241569
Rin97_41 in97_40 in97_41 9.241569
Rin97_42 in97_41 in97_42 9.241569
Rin97_43 in97_42 in97_43 9.241569
Rin97_44 in97_43 in97_44 9.241569
Rin97_45 in97_44 in97_45 9.241569
Rin97_46 in97_45 in97_46 9.241569
Rin97_47 in97_46 in97_47 9.241569
Rin97_48 in97_47 in97_48 9.241569
Rin97_49 in97_48 in97_49 9.241569
Rin97_50 in97_49 in97_50 9.241569
Rin97_51 in97_50 in97_51 9.241569
Rin97_52 in97_51 in97_52 9.241569
Rin97_53 in97_52 in97_53 9.241569
Rin97_54 in97_53 in97_54 9.241569
Rin97_55 in97_54 in97_55 9.241569
Rin97_56 in97_55 in97_56 9.241569
Rin97_57 in97 in97_57 9.241569
Rin97_58 in97_57 in97_58 9.241569
Rin97_59 in97_58 in97_59 9.241569
Rin97_60 in97_59 in97_60 9.241569
Rin97_61 in97_60 in97_61 9.241569
Rin97_62 in97_61 in97_62 9.241569
Rin97_63 in97_62 in97_63 9.241569
Rin97_64 in97_63 in97_64 9.241569
Rin97_65 in97_64 in97_65 9.241569
Rin97_66 in97_65 in97_66 9.241569
Rin97_67 in97_66 in97_67 9.241569
Rin97_68 in97_67 in97_68 9.241569
Rin97_69 in97_68 in97_69 9.241569
Rin97_70 in97_69 in97_70 9.241569
Rin97_71 in97_70 in97_71 9.241569
Rin97_72 in97_71 in97_72 9.241569
Rin97_73 in97_72 in97_73 9.241569
Rin97_74 in97_73 in97_74 9.241569
Rin97_75 in97_74 in97_75 9.241569
Rin97_76 in97_75 in97_76 9.241569
Rin97_77 in97_76 in97_77 9.241569
Rin97_78 in97_77 in97_78 9.241569
Rin97_79 in97_78 in97_79 9.241569
Rin97_80 in97_79 in97_80 9.241569
Rin97_81 in97_80 in97_81 9.241569
Rin97_82 in97_81 in97_82 9.241569
Rin97_83 in97_82 in97_83 9.241569
Rin97_84 in97_83 in97_84 9.241569
Rin98_1 in98 in98_1 9.241569
Rin98_2 in98_1 in98_2 9.241569
Rin98_3 in98_2 in98_3 9.241569
Rin98_4 in98_3 in98_4 9.241569
Rin98_5 in98_4 in98_5 9.241569
Rin98_6 in98_5 in98_6 9.241569
Rin98_7 in98_6 in98_7 9.241569
Rin98_8 in98_7 in98_8 9.241569
Rin98_9 in98_8 in98_9 9.241569
Rin98_10 in98_9 in98_10 9.241569
Rin98_11 in98_10 in98_11 9.241569
Rin98_12 in98_11 in98_12 9.241569
Rin98_13 in98_12 in98_13 9.241569
Rin98_14 in98_13 in98_14 9.241569
Rin98_15 in98_14 in98_15 9.241569
Rin98_16 in98_15 in98_16 9.241569
Rin98_17 in98_16 in98_17 9.241569
Rin98_18 in98_17 in98_18 9.241569
Rin98_19 in98_18 in98_19 9.241569
Rin98_20 in98_19 in98_20 9.241569
Rin98_21 in98_20 in98_21 9.241569
Rin98_22 in98_21 in98_22 9.241569
Rin98_23 in98_22 in98_23 9.241569
Rin98_24 in98_23 in98_24 9.241569
Rin98_25 in98_24 in98_25 9.241569
Rin98_26 in98_25 in98_26 9.241569
Rin98_27 in98_26 in98_27 9.241569
Rin98_28 in98_27 in98_28 9.241569
Rin98_29 in98 in98_29 9.241569
Rin98_30 in98_29 in98_30 9.241569
Rin98_31 in98_30 in98_31 9.241569
Rin98_32 in98_31 in98_32 9.241569
Rin98_33 in98_32 in98_33 9.241569
Rin98_34 in98_33 in98_34 9.241569
Rin98_35 in98_34 in98_35 9.241569
Rin98_36 in98_35 in98_36 9.241569
Rin98_37 in98_36 in98_37 9.241569
Rin98_38 in98_37 in98_38 9.241569
Rin98_39 in98_38 in98_39 9.241569
Rin98_40 in98_39 in98_40 9.241569
Rin98_41 in98_40 in98_41 9.241569
Rin98_42 in98_41 in98_42 9.241569
Rin98_43 in98_42 in98_43 9.241569
Rin98_44 in98_43 in98_44 9.241569
Rin98_45 in98_44 in98_45 9.241569
Rin98_46 in98_45 in98_46 9.241569
Rin98_47 in98_46 in98_47 9.241569
Rin98_48 in98_47 in98_48 9.241569
Rin98_49 in98_48 in98_49 9.241569
Rin98_50 in98_49 in98_50 9.241569
Rin98_51 in98_50 in98_51 9.241569
Rin98_52 in98_51 in98_52 9.241569
Rin98_53 in98_52 in98_53 9.241569
Rin98_54 in98_53 in98_54 9.241569
Rin98_55 in98_54 in98_55 9.241569
Rin98_56 in98_55 in98_56 9.241569
Rin98_57 in98 in98_57 9.241569
Rin98_58 in98_57 in98_58 9.241569
Rin98_59 in98_58 in98_59 9.241569
Rin98_60 in98_59 in98_60 9.241569
Rin98_61 in98_60 in98_61 9.241569
Rin98_62 in98_61 in98_62 9.241569
Rin98_63 in98_62 in98_63 9.241569
Rin98_64 in98_63 in98_64 9.241569
Rin98_65 in98_64 in98_65 9.241569
Rin98_66 in98_65 in98_66 9.241569
Rin98_67 in98_66 in98_67 9.241569
Rin98_68 in98_67 in98_68 9.241569
Rin98_69 in98_68 in98_69 9.241569
Rin98_70 in98_69 in98_70 9.241569
Rin98_71 in98_70 in98_71 9.241569
Rin98_72 in98_71 in98_72 9.241569
Rin98_73 in98_72 in98_73 9.241569
Rin98_74 in98_73 in98_74 9.241569
Rin98_75 in98_74 in98_75 9.241569
Rin98_76 in98_75 in98_76 9.241569
Rin98_77 in98_76 in98_77 9.241569
Rin98_78 in98_77 in98_78 9.241569
Rin98_79 in98_78 in98_79 9.241569
Rin98_80 in98_79 in98_80 9.241569
Rin98_81 in98_80 in98_81 9.241569
Rin98_82 in98_81 in98_82 9.241569
Rin98_83 in98_82 in98_83 9.241569
Rin98_84 in98_83 in98_84 9.241569
Rin99_1 in99 in99_1 9.241569
Rin99_2 in99_1 in99_2 9.241569
Rin99_3 in99_2 in99_3 9.241569
Rin99_4 in99_3 in99_4 9.241569
Rin99_5 in99_4 in99_5 9.241569
Rin99_6 in99_5 in99_6 9.241569
Rin99_7 in99_6 in99_7 9.241569
Rin99_8 in99_7 in99_8 9.241569
Rin99_9 in99_8 in99_9 9.241569
Rin99_10 in99_9 in99_10 9.241569
Rin99_11 in99_10 in99_11 9.241569
Rin99_12 in99_11 in99_12 9.241569
Rin99_13 in99_12 in99_13 9.241569
Rin99_14 in99_13 in99_14 9.241569
Rin99_15 in99_14 in99_15 9.241569
Rin99_16 in99_15 in99_16 9.241569
Rin99_17 in99_16 in99_17 9.241569
Rin99_18 in99_17 in99_18 9.241569
Rin99_19 in99_18 in99_19 9.241569
Rin99_20 in99_19 in99_20 9.241569
Rin99_21 in99_20 in99_21 9.241569
Rin99_22 in99_21 in99_22 9.241569
Rin99_23 in99_22 in99_23 9.241569
Rin99_24 in99_23 in99_24 9.241569
Rin99_25 in99_24 in99_25 9.241569
Rin99_26 in99_25 in99_26 9.241569
Rin99_27 in99_26 in99_27 9.241569
Rin99_28 in99_27 in99_28 9.241569
Rin99_29 in99 in99_29 9.241569
Rin99_30 in99_29 in99_30 9.241569
Rin99_31 in99_30 in99_31 9.241569
Rin99_32 in99_31 in99_32 9.241569
Rin99_33 in99_32 in99_33 9.241569
Rin99_34 in99_33 in99_34 9.241569
Rin99_35 in99_34 in99_35 9.241569
Rin99_36 in99_35 in99_36 9.241569
Rin99_37 in99_36 in99_37 9.241569
Rin99_38 in99_37 in99_38 9.241569
Rin99_39 in99_38 in99_39 9.241569
Rin99_40 in99_39 in99_40 9.241569
Rin99_41 in99_40 in99_41 9.241569
Rin99_42 in99_41 in99_42 9.241569
Rin99_43 in99_42 in99_43 9.241569
Rin99_44 in99_43 in99_44 9.241569
Rin99_45 in99_44 in99_45 9.241569
Rin99_46 in99_45 in99_46 9.241569
Rin99_47 in99_46 in99_47 9.241569
Rin99_48 in99_47 in99_48 9.241569
Rin99_49 in99_48 in99_49 9.241569
Rin99_50 in99_49 in99_50 9.241569
Rin99_51 in99_50 in99_51 9.241569
Rin99_52 in99_51 in99_52 9.241569
Rin99_53 in99_52 in99_53 9.241569
Rin99_54 in99_53 in99_54 9.241569
Rin99_55 in99_54 in99_55 9.241569
Rin99_56 in99_55 in99_56 9.241569
Rin99_57 in99 in99_57 9.241569
Rin99_58 in99_57 in99_58 9.241569
Rin99_59 in99_58 in99_59 9.241569
Rin99_60 in99_59 in99_60 9.241569
Rin99_61 in99_60 in99_61 9.241569
Rin99_62 in99_61 in99_62 9.241569
Rin99_63 in99_62 in99_63 9.241569
Rin99_64 in99_63 in99_64 9.241569
Rin99_65 in99_64 in99_65 9.241569
Rin99_66 in99_65 in99_66 9.241569
Rin99_67 in99_66 in99_67 9.241569
Rin99_68 in99_67 in99_68 9.241569
Rin99_69 in99_68 in99_69 9.241569
Rin99_70 in99_69 in99_70 9.241569
Rin99_71 in99_70 in99_71 9.241569
Rin99_72 in99_71 in99_72 9.241569
Rin99_73 in99_72 in99_73 9.241569
Rin99_74 in99_73 in99_74 9.241569
Rin99_75 in99_74 in99_75 9.241569
Rin99_76 in99_75 in99_76 9.241569
Rin99_77 in99_76 in99_77 9.241569
Rin99_78 in99_77 in99_78 9.241569
Rin99_79 in99_78 in99_79 9.241569
Rin99_80 in99_79 in99_80 9.241569
Rin99_81 in99_80 in99_81 9.241569
Rin99_82 in99_81 in99_82 9.241569
Rin99_83 in99_82 in99_83 9.241569
Rin99_84 in99_83 in99_84 9.241569
Rin100_1 in100 in100_1 9.241569
Rin100_2 in100_1 in100_2 9.241569
Rin100_3 in100_2 in100_3 9.241569
Rin100_4 in100_3 in100_4 9.241569
Rin100_5 in100_4 in100_5 9.241569
Rin100_6 in100_5 in100_6 9.241569
Rin100_7 in100_6 in100_7 9.241569
Rin100_8 in100_7 in100_8 9.241569
Rin100_9 in100_8 in100_9 9.241569
Rin100_10 in100_9 in100_10 9.241569
Rin100_11 in100_10 in100_11 9.241569
Rin100_12 in100_11 in100_12 9.241569
Rin100_13 in100_12 in100_13 9.241569
Rin100_14 in100_13 in100_14 9.241569
Rin100_15 in100_14 in100_15 9.241569
Rin100_16 in100_15 in100_16 9.241569
Rin100_17 in100_16 in100_17 9.241569
Rin100_18 in100_17 in100_18 9.241569
Rin100_19 in100_18 in100_19 9.241569
Rin100_20 in100_19 in100_20 9.241569
Rin100_21 in100_20 in100_21 9.241569
Rin100_22 in100_21 in100_22 9.241569
Rin100_23 in100_22 in100_23 9.241569
Rin100_24 in100_23 in100_24 9.241569
Rin100_25 in100_24 in100_25 9.241569
Rin100_26 in100_25 in100_26 9.241569
Rin100_27 in100_26 in100_27 9.241569
Rin100_28 in100_27 in100_28 9.241569
Rin100_29 in100 in100_29 9.241569
Rin100_30 in100_29 in100_30 9.241569
Rin100_31 in100_30 in100_31 9.241569
Rin100_32 in100_31 in100_32 9.241569
Rin100_33 in100_32 in100_33 9.241569
Rin100_34 in100_33 in100_34 9.241569
Rin100_35 in100_34 in100_35 9.241569
Rin100_36 in100_35 in100_36 9.241569
Rin100_37 in100_36 in100_37 9.241569
Rin100_38 in100_37 in100_38 9.241569
Rin100_39 in100_38 in100_39 9.241569
Rin100_40 in100_39 in100_40 9.241569
Rin100_41 in100_40 in100_41 9.241569
Rin100_42 in100_41 in100_42 9.241569
Rin100_43 in100_42 in100_43 9.241569
Rin100_44 in100_43 in100_44 9.241569
Rin100_45 in100_44 in100_45 9.241569
Rin100_46 in100_45 in100_46 9.241569
Rin100_47 in100_46 in100_47 9.241569
Rin100_48 in100_47 in100_48 9.241569
Rin100_49 in100_48 in100_49 9.241569
Rin100_50 in100_49 in100_50 9.241569
Rin100_51 in100_50 in100_51 9.241569
Rin100_52 in100_51 in100_52 9.241569
Rin100_53 in100_52 in100_53 9.241569
Rin100_54 in100_53 in100_54 9.241569
Rin100_55 in100_54 in100_55 9.241569
Rin100_56 in100_55 in100_56 9.241569
Rin100_57 in100 in100_57 9.241569
Rin100_58 in100_57 in100_58 9.241569
Rin100_59 in100_58 in100_59 9.241569
Rin100_60 in100_59 in100_60 9.241569
Rin100_61 in100_60 in100_61 9.241569
Rin100_62 in100_61 in100_62 9.241569
Rin100_63 in100_62 in100_63 9.241569
Rin100_64 in100_63 in100_64 9.241569
Rin100_65 in100_64 in100_65 9.241569
Rin100_66 in100_65 in100_66 9.241569
Rin100_67 in100_66 in100_67 9.241569
Rin100_68 in100_67 in100_68 9.241569
Rin100_69 in100_68 in100_69 9.241569
Rin100_70 in100_69 in100_70 9.241569
Rin100_71 in100_70 in100_71 9.241569
Rin100_72 in100_71 in100_72 9.241569
Rin100_73 in100_72 in100_73 9.241569
Rin100_74 in100_73 in100_74 9.241569
Rin100_75 in100_74 in100_75 9.241569
Rin100_76 in100_75 in100_76 9.241569
Rin100_77 in100_76 in100_77 9.241569
Rin100_78 in100_77 in100_78 9.241569
Rin100_79 in100_78 in100_79 9.241569
Rin100_80 in100_79 in100_80 9.241569
Rin100_81 in100_80 in100_81 9.241569
Rin100_82 in100_81 in100_82 9.241569
Rin100_83 in100_82 in100_83 9.241569
Rin100_84 in100_83 in100_84 9.241569
Rin101_1 in101 in101_1 9.241569
Rin101_2 in101_1 in101_2 9.241569
Rin101_3 in101_2 in101_3 9.241569
Rin101_4 in101_3 in101_4 9.241569
Rin101_5 in101_4 in101_5 9.241569
Rin101_6 in101_5 in101_6 9.241569
Rin101_7 in101_6 in101_7 9.241569
Rin101_8 in101_7 in101_8 9.241569
Rin101_9 in101_8 in101_9 9.241569
Rin101_10 in101_9 in101_10 9.241569
Rin101_11 in101_10 in101_11 9.241569
Rin101_12 in101_11 in101_12 9.241569
Rin101_13 in101_12 in101_13 9.241569
Rin101_14 in101_13 in101_14 9.241569
Rin101_15 in101_14 in101_15 9.241569
Rin101_16 in101_15 in101_16 9.241569
Rin101_17 in101_16 in101_17 9.241569
Rin101_18 in101_17 in101_18 9.241569
Rin101_19 in101_18 in101_19 9.241569
Rin101_20 in101_19 in101_20 9.241569
Rin101_21 in101_20 in101_21 9.241569
Rin101_22 in101_21 in101_22 9.241569
Rin101_23 in101_22 in101_23 9.241569
Rin101_24 in101_23 in101_24 9.241569
Rin101_25 in101_24 in101_25 9.241569
Rin101_26 in101_25 in101_26 9.241569
Rin101_27 in101_26 in101_27 9.241569
Rin101_28 in101_27 in101_28 9.241569
Rin101_29 in101 in101_29 9.241569
Rin101_30 in101_29 in101_30 9.241569
Rin101_31 in101_30 in101_31 9.241569
Rin101_32 in101_31 in101_32 9.241569
Rin101_33 in101_32 in101_33 9.241569
Rin101_34 in101_33 in101_34 9.241569
Rin101_35 in101_34 in101_35 9.241569
Rin101_36 in101_35 in101_36 9.241569
Rin101_37 in101_36 in101_37 9.241569
Rin101_38 in101_37 in101_38 9.241569
Rin101_39 in101_38 in101_39 9.241569
Rin101_40 in101_39 in101_40 9.241569
Rin101_41 in101_40 in101_41 9.241569
Rin101_42 in101_41 in101_42 9.241569
Rin101_43 in101_42 in101_43 9.241569
Rin101_44 in101_43 in101_44 9.241569
Rin101_45 in101_44 in101_45 9.241569
Rin101_46 in101_45 in101_46 9.241569
Rin101_47 in101_46 in101_47 9.241569
Rin101_48 in101_47 in101_48 9.241569
Rin101_49 in101_48 in101_49 9.241569
Rin101_50 in101_49 in101_50 9.241569
Rin101_51 in101_50 in101_51 9.241569
Rin101_52 in101_51 in101_52 9.241569
Rin101_53 in101_52 in101_53 9.241569
Rin101_54 in101_53 in101_54 9.241569
Rin101_55 in101_54 in101_55 9.241569
Rin101_56 in101_55 in101_56 9.241569
Rin101_57 in101 in101_57 9.241569
Rin101_58 in101_57 in101_58 9.241569
Rin101_59 in101_58 in101_59 9.241569
Rin101_60 in101_59 in101_60 9.241569
Rin101_61 in101_60 in101_61 9.241569
Rin101_62 in101_61 in101_62 9.241569
Rin101_63 in101_62 in101_63 9.241569
Rin101_64 in101_63 in101_64 9.241569
Rin101_65 in101_64 in101_65 9.241569
Rin101_66 in101_65 in101_66 9.241569
Rin101_67 in101_66 in101_67 9.241569
Rin101_68 in101_67 in101_68 9.241569
Rin101_69 in101_68 in101_69 9.241569
Rin101_70 in101_69 in101_70 9.241569
Rin101_71 in101_70 in101_71 9.241569
Rin101_72 in101_71 in101_72 9.241569
Rin101_73 in101_72 in101_73 9.241569
Rin101_74 in101_73 in101_74 9.241569
Rin101_75 in101_74 in101_75 9.241569
Rin101_76 in101_75 in101_76 9.241569
Rin101_77 in101_76 in101_77 9.241569
Rin101_78 in101_77 in101_78 9.241569
Rin101_79 in101_78 in101_79 9.241569
Rin101_80 in101_79 in101_80 9.241569
Rin101_81 in101_80 in101_81 9.241569
Rin101_82 in101_81 in101_82 9.241569
Rin101_83 in101_82 in101_83 9.241569
Rin101_84 in101_83 in101_84 9.241569
Rin102_1 in102 in102_1 9.241569
Rin102_2 in102_1 in102_2 9.241569
Rin102_3 in102_2 in102_3 9.241569
Rin102_4 in102_3 in102_4 9.241569
Rin102_5 in102_4 in102_5 9.241569
Rin102_6 in102_5 in102_6 9.241569
Rin102_7 in102_6 in102_7 9.241569
Rin102_8 in102_7 in102_8 9.241569
Rin102_9 in102_8 in102_9 9.241569
Rin102_10 in102_9 in102_10 9.241569
Rin102_11 in102_10 in102_11 9.241569
Rin102_12 in102_11 in102_12 9.241569
Rin102_13 in102_12 in102_13 9.241569
Rin102_14 in102_13 in102_14 9.241569
Rin102_15 in102_14 in102_15 9.241569
Rin102_16 in102_15 in102_16 9.241569
Rin102_17 in102_16 in102_17 9.241569
Rin102_18 in102_17 in102_18 9.241569
Rin102_19 in102_18 in102_19 9.241569
Rin102_20 in102_19 in102_20 9.241569
Rin102_21 in102_20 in102_21 9.241569
Rin102_22 in102_21 in102_22 9.241569
Rin102_23 in102_22 in102_23 9.241569
Rin102_24 in102_23 in102_24 9.241569
Rin102_25 in102_24 in102_25 9.241569
Rin102_26 in102_25 in102_26 9.241569
Rin102_27 in102_26 in102_27 9.241569
Rin102_28 in102_27 in102_28 9.241569
Rin102_29 in102 in102_29 9.241569
Rin102_30 in102_29 in102_30 9.241569
Rin102_31 in102_30 in102_31 9.241569
Rin102_32 in102_31 in102_32 9.241569
Rin102_33 in102_32 in102_33 9.241569
Rin102_34 in102_33 in102_34 9.241569
Rin102_35 in102_34 in102_35 9.241569
Rin102_36 in102_35 in102_36 9.241569
Rin102_37 in102_36 in102_37 9.241569
Rin102_38 in102_37 in102_38 9.241569
Rin102_39 in102_38 in102_39 9.241569
Rin102_40 in102_39 in102_40 9.241569
Rin102_41 in102_40 in102_41 9.241569
Rin102_42 in102_41 in102_42 9.241569
Rin102_43 in102_42 in102_43 9.241569
Rin102_44 in102_43 in102_44 9.241569
Rin102_45 in102_44 in102_45 9.241569
Rin102_46 in102_45 in102_46 9.241569
Rin102_47 in102_46 in102_47 9.241569
Rin102_48 in102_47 in102_48 9.241569
Rin102_49 in102_48 in102_49 9.241569
Rin102_50 in102_49 in102_50 9.241569
Rin102_51 in102_50 in102_51 9.241569
Rin102_52 in102_51 in102_52 9.241569
Rin102_53 in102_52 in102_53 9.241569
Rin102_54 in102_53 in102_54 9.241569
Rin102_55 in102_54 in102_55 9.241569
Rin102_56 in102_55 in102_56 9.241569
Rin102_57 in102 in102_57 9.241569
Rin102_58 in102_57 in102_58 9.241569
Rin102_59 in102_58 in102_59 9.241569
Rin102_60 in102_59 in102_60 9.241569
Rin102_61 in102_60 in102_61 9.241569
Rin102_62 in102_61 in102_62 9.241569
Rin102_63 in102_62 in102_63 9.241569
Rin102_64 in102_63 in102_64 9.241569
Rin102_65 in102_64 in102_65 9.241569
Rin102_66 in102_65 in102_66 9.241569
Rin102_67 in102_66 in102_67 9.241569
Rin102_68 in102_67 in102_68 9.241569
Rin102_69 in102_68 in102_69 9.241569
Rin102_70 in102_69 in102_70 9.241569
Rin102_71 in102_70 in102_71 9.241569
Rin102_72 in102_71 in102_72 9.241569
Rin102_73 in102_72 in102_73 9.241569
Rin102_74 in102_73 in102_74 9.241569
Rin102_75 in102_74 in102_75 9.241569
Rin102_76 in102_75 in102_76 9.241569
Rin102_77 in102_76 in102_77 9.241569
Rin102_78 in102_77 in102_78 9.241569
Rin102_79 in102_78 in102_79 9.241569
Rin102_80 in102_79 in102_80 9.241569
Rin102_81 in102_80 in102_81 9.241569
Rin102_82 in102_81 in102_82 9.241569
Rin102_83 in102_82 in102_83 9.241569
Rin102_84 in102_83 in102_84 9.241569
Rin103_1 in103 in103_1 9.241569
Rin103_2 in103_1 in103_2 9.241569
Rin103_3 in103_2 in103_3 9.241569
Rin103_4 in103_3 in103_4 9.241569
Rin103_5 in103_4 in103_5 9.241569
Rin103_6 in103_5 in103_6 9.241569
Rin103_7 in103_6 in103_7 9.241569
Rin103_8 in103_7 in103_8 9.241569
Rin103_9 in103_8 in103_9 9.241569
Rin103_10 in103_9 in103_10 9.241569
Rin103_11 in103_10 in103_11 9.241569
Rin103_12 in103_11 in103_12 9.241569
Rin103_13 in103_12 in103_13 9.241569
Rin103_14 in103_13 in103_14 9.241569
Rin103_15 in103_14 in103_15 9.241569
Rin103_16 in103_15 in103_16 9.241569
Rin103_17 in103_16 in103_17 9.241569
Rin103_18 in103_17 in103_18 9.241569
Rin103_19 in103_18 in103_19 9.241569
Rin103_20 in103_19 in103_20 9.241569
Rin103_21 in103_20 in103_21 9.241569
Rin103_22 in103_21 in103_22 9.241569
Rin103_23 in103_22 in103_23 9.241569
Rin103_24 in103_23 in103_24 9.241569
Rin103_25 in103_24 in103_25 9.241569
Rin103_26 in103_25 in103_26 9.241569
Rin103_27 in103_26 in103_27 9.241569
Rin103_28 in103_27 in103_28 9.241569
Rin103_29 in103 in103_29 9.241569
Rin103_30 in103_29 in103_30 9.241569
Rin103_31 in103_30 in103_31 9.241569
Rin103_32 in103_31 in103_32 9.241569
Rin103_33 in103_32 in103_33 9.241569
Rin103_34 in103_33 in103_34 9.241569
Rin103_35 in103_34 in103_35 9.241569
Rin103_36 in103_35 in103_36 9.241569
Rin103_37 in103_36 in103_37 9.241569
Rin103_38 in103_37 in103_38 9.241569
Rin103_39 in103_38 in103_39 9.241569
Rin103_40 in103_39 in103_40 9.241569
Rin103_41 in103_40 in103_41 9.241569
Rin103_42 in103_41 in103_42 9.241569
Rin103_43 in103_42 in103_43 9.241569
Rin103_44 in103_43 in103_44 9.241569
Rin103_45 in103_44 in103_45 9.241569
Rin103_46 in103_45 in103_46 9.241569
Rin103_47 in103_46 in103_47 9.241569
Rin103_48 in103_47 in103_48 9.241569
Rin103_49 in103_48 in103_49 9.241569
Rin103_50 in103_49 in103_50 9.241569
Rin103_51 in103_50 in103_51 9.241569
Rin103_52 in103_51 in103_52 9.241569
Rin103_53 in103_52 in103_53 9.241569
Rin103_54 in103_53 in103_54 9.241569
Rin103_55 in103_54 in103_55 9.241569
Rin103_56 in103_55 in103_56 9.241569
Rin103_57 in103 in103_57 9.241569
Rin103_58 in103_57 in103_58 9.241569
Rin103_59 in103_58 in103_59 9.241569
Rin103_60 in103_59 in103_60 9.241569
Rin103_61 in103_60 in103_61 9.241569
Rin103_62 in103_61 in103_62 9.241569
Rin103_63 in103_62 in103_63 9.241569
Rin103_64 in103_63 in103_64 9.241569
Rin103_65 in103_64 in103_65 9.241569
Rin103_66 in103_65 in103_66 9.241569
Rin103_67 in103_66 in103_67 9.241569
Rin103_68 in103_67 in103_68 9.241569
Rin103_69 in103_68 in103_69 9.241569
Rin103_70 in103_69 in103_70 9.241569
Rin103_71 in103_70 in103_71 9.241569
Rin103_72 in103_71 in103_72 9.241569
Rin103_73 in103_72 in103_73 9.241569
Rin103_74 in103_73 in103_74 9.241569
Rin103_75 in103_74 in103_75 9.241569
Rin103_76 in103_75 in103_76 9.241569
Rin103_77 in103_76 in103_77 9.241569
Rin103_78 in103_77 in103_78 9.241569
Rin103_79 in103_78 in103_79 9.241569
Rin103_80 in103_79 in103_80 9.241569
Rin103_81 in103_80 in103_81 9.241569
Rin103_82 in103_81 in103_82 9.241569
Rin103_83 in103_82 in103_83 9.241569
Rin103_84 in103_83 in103_84 9.241569
Rin104_1 in104 in104_1 9.241569
Rin104_2 in104_1 in104_2 9.241569
Rin104_3 in104_2 in104_3 9.241569
Rin104_4 in104_3 in104_4 9.241569
Rin104_5 in104_4 in104_5 9.241569
Rin104_6 in104_5 in104_6 9.241569
Rin104_7 in104_6 in104_7 9.241569
Rin104_8 in104_7 in104_8 9.241569
Rin104_9 in104_8 in104_9 9.241569
Rin104_10 in104_9 in104_10 9.241569
Rin104_11 in104_10 in104_11 9.241569
Rin104_12 in104_11 in104_12 9.241569
Rin104_13 in104_12 in104_13 9.241569
Rin104_14 in104_13 in104_14 9.241569
Rin104_15 in104_14 in104_15 9.241569
Rin104_16 in104_15 in104_16 9.241569
Rin104_17 in104_16 in104_17 9.241569
Rin104_18 in104_17 in104_18 9.241569
Rin104_19 in104_18 in104_19 9.241569
Rin104_20 in104_19 in104_20 9.241569
Rin104_21 in104_20 in104_21 9.241569
Rin104_22 in104_21 in104_22 9.241569
Rin104_23 in104_22 in104_23 9.241569
Rin104_24 in104_23 in104_24 9.241569
Rin104_25 in104_24 in104_25 9.241569
Rin104_26 in104_25 in104_26 9.241569
Rin104_27 in104_26 in104_27 9.241569
Rin104_28 in104_27 in104_28 9.241569
Rin104_29 in104 in104_29 9.241569
Rin104_30 in104_29 in104_30 9.241569
Rin104_31 in104_30 in104_31 9.241569
Rin104_32 in104_31 in104_32 9.241569
Rin104_33 in104_32 in104_33 9.241569
Rin104_34 in104_33 in104_34 9.241569
Rin104_35 in104_34 in104_35 9.241569
Rin104_36 in104_35 in104_36 9.241569
Rin104_37 in104_36 in104_37 9.241569
Rin104_38 in104_37 in104_38 9.241569
Rin104_39 in104_38 in104_39 9.241569
Rin104_40 in104_39 in104_40 9.241569
Rin104_41 in104_40 in104_41 9.241569
Rin104_42 in104_41 in104_42 9.241569
Rin104_43 in104_42 in104_43 9.241569
Rin104_44 in104_43 in104_44 9.241569
Rin104_45 in104_44 in104_45 9.241569
Rin104_46 in104_45 in104_46 9.241569
Rin104_47 in104_46 in104_47 9.241569
Rin104_48 in104_47 in104_48 9.241569
Rin104_49 in104_48 in104_49 9.241569
Rin104_50 in104_49 in104_50 9.241569
Rin104_51 in104_50 in104_51 9.241569
Rin104_52 in104_51 in104_52 9.241569
Rin104_53 in104_52 in104_53 9.241569
Rin104_54 in104_53 in104_54 9.241569
Rin104_55 in104_54 in104_55 9.241569
Rin104_56 in104_55 in104_56 9.241569
Rin104_57 in104 in104_57 9.241569
Rin104_58 in104_57 in104_58 9.241569
Rin104_59 in104_58 in104_59 9.241569
Rin104_60 in104_59 in104_60 9.241569
Rin104_61 in104_60 in104_61 9.241569
Rin104_62 in104_61 in104_62 9.241569
Rin104_63 in104_62 in104_63 9.241569
Rin104_64 in104_63 in104_64 9.241569
Rin104_65 in104_64 in104_65 9.241569
Rin104_66 in104_65 in104_66 9.241569
Rin104_67 in104_66 in104_67 9.241569
Rin104_68 in104_67 in104_68 9.241569
Rin104_69 in104_68 in104_69 9.241569
Rin104_70 in104_69 in104_70 9.241569
Rin104_71 in104_70 in104_71 9.241569
Rin104_72 in104_71 in104_72 9.241569
Rin104_73 in104_72 in104_73 9.241569
Rin104_74 in104_73 in104_74 9.241569
Rin104_75 in104_74 in104_75 9.241569
Rin104_76 in104_75 in104_76 9.241569
Rin104_77 in104_76 in104_77 9.241569
Rin104_78 in104_77 in104_78 9.241569
Rin104_79 in104_78 in104_79 9.241569
Rin104_80 in104_79 in104_80 9.241569
Rin104_81 in104_80 in104_81 9.241569
Rin104_82 in104_81 in104_82 9.241569
Rin104_83 in104_82 in104_83 9.241569
Rin104_84 in104_83 in104_84 9.241569
Rin105_1 in105 in105_1 9.241569
Rin105_2 in105_1 in105_2 9.241569
Rin105_3 in105_2 in105_3 9.241569
Rin105_4 in105_3 in105_4 9.241569
Rin105_5 in105_4 in105_5 9.241569
Rin105_6 in105_5 in105_6 9.241569
Rin105_7 in105_6 in105_7 9.241569
Rin105_8 in105_7 in105_8 9.241569
Rin105_9 in105_8 in105_9 9.241569
Rin105_10 in105_9 in105_10 9.241569
Rin105_11 in105_10 in105_11 9.241569
Rin105_12 in105_11 in105_12 9.241569
Rin105_13 in105_12 in105_13 9.241569
Rin105_14 in105_13 in105_14 9.241569
Rin105_15 in105_14 in105_15 9.241569
Rin105_16 in105_15 in105_16 9.241569
Rin105_17 in105_16 in105_17 9.241569
Rin105_18 in105_17 in105_18 9.241569
Rin105_19 in105_18 in105_19 9.241569
Rin105_20 in105_19 in105_20 9.241569
Rin105_21 in105_20 in105_21 9.241569
Rin105_22 in105_21 in105_22 9.241569
Rin105_23 in105_22 in105_23 9.241569
Rin105_24 in105_23 in105_24 9.241569
Rin105_25 in105_24 in105_25 9.241569
Rin105_26 in105_25 in105_26 9.241569
Rin105_27 in105_26 in105_27 9.241569
Rin105_28 in105_27 in105_28 9.241569
Rin105_29 in105 in105_29 9.241569
Rin105_30 in105_29 in105_30 9.241569
Rin105_31 in105_30 in105_31 9.241569
Rin105_32 in105_31 in105_32 9.241569
Rin105_33 in105_32 in105_33 9.241569
Rin105_34 in105_33 in105_34 9.241569
Rin105_35 in105_34 in105_35 9.241569
Rin105_36 in105_35 in105_36 9.241569
Rin105_37 in105_36 in105_37 9.241569
Rin105_38 in105_37 in105_38 9.241569
Rin105_39 in105_38 in105_39 9.241569
Rin105_40 in105_39 in105_40 9.241569
Rin105_41 in105_40 in105_41 9.241569
Rin105_42 in105_41 in105_42 9.241569
Rin105_43 in105_42 in105_43 9.241569
Rin105_44 in105_43 in105_44 9.241569
Rin105_45 in105_44 in105_45 9.241569
Rin105_46 in105_45 in105_46 9.241569
Rin105_47 in105_46 in105_47 9.241569
Rin105_48 in105_47 in105_48 9.241569
Rin105_49 in105_48 in105_49 9.241569
Rin105_50 in105_49 in105_50 9.241569
Rin105_51 in105_50 in105_51 9.241569
Rin105_52 in105_51 in105_52 9.241569
Rin105_53 in105_52 in105_53 9.241569
Rin105_54 in105_53 in105_54 9.241569
Rin105_55 in105_54 in105_55 9.241569
Rin105_56 in105_55 in105_56 9.241569
Rin105_57 in105 in105_57 9.241569
Rin105_58 in105_57 in105_58 9.241569
Rin105_59 in105_58 in105_59 9.241569
Rin105_60 in105_59 in105_60 9.241569
Rin105_61 in105_60 in105_61 9.241569
Rin105_62 in105_61 in105_62 9.241569
Rin105_63 in105_62 in105_63 9.241569
Rin105_64 in105_63 in105_64 9.241569
Rin105_65 in105_64 in105_65 9.241569
Rin105_66 in105_65 in105_66 9.241569
Rin105_67 in105_66 in105_67 9.241569
Rin105_68 in105_67 in105_68 9.241569
Rin105_69 in105_68 in105_69 9.241569
Rin105_70 in105_69 in105_70 9.241569
Rin105_71 in105_70 in105_71 9.241569
Rin105_72 in105_71 in105_72 9.241569
Rin105_73 in105_72 in105_73 9.241569
Rin105_74 in105_73 in105_74 9.241569
Rin105_75 in105_74 in105_75 9.241569
Rin105_76 in105_75 in105_76 9.241569
Rin105_77 in105_76 in105_77 9.241569
Rin105_78 in105_77 in105_78 9.241569
Rin105_79 in105_78 in105_79 9.241569
Rin105_80 in105_79 in105_80 9.241569
Rin105_81 in105_80 in105_81 9.241569
Rin105_82 in105_81 in105_82 9.241569
Rin105_83 in105_82 in105_83 9.241569
Rin105_84 in105_83 in105_84 9.241569
Rin106_1 in106 in106_1 9.241569
Rin106_2 in106_1 in106_2 9.241569
Rin106_3 in106_2 in106_3 9.241569
Rin106_4 in106_3 in106_4 9.241569
Rin106_5 in106_4 in106_5 9.241569
Rin106_6 in106_5 in106_6 9.241569
Rin106_7 in106_6 in106_7 9.241569
Rin106_8 in106_7 in106_8 9.241569
Rin106_9 in106_8 in106_9 9.241569
Rin106_10 in106_9 in106_10 9.241569
Rin106_11 in106_10 in106_11 9.241569
Rin106_12 in106_11 in106_12 9.241569
Rin106_13 in106_12 in106_13 9.241569
Rin106_14 in106_13 in106_14 9.241569
Rin106_15 in106_14 in106_15 9.241569
Rin106_16 in106_15 in106_16 9.241569
Rin106_17 in106_16 in106_17 9.241569
Rin106_18 in106_17 in106_18 9.241569
Rin106_19 in106_18 in106_19 9.241569
Rin106_20 in106_19 in106_20 9.241569
Rin106_21 in106_20 in106_21 9.241569
Rin106_22 in106_21 in106_22 9.241569
Rin106_23 in106_22 in106_23 9.241569
Rin106_24 in106_23 in106_24 9.241569
Rin106_25 in106_24 in106_25 9.241569
Rin106_26 in106_25 in106_26 9.241569
Rin106_27 in106_26 in106_27 9.241569
Rin106_28 in106_27 in106_28 9.241569
Rin106_29 in106 in106_29 9.241569
Rin106_30 in106_29 in106_30 9.241569
Rin106_31 in106_30 in106_31 9.241569
Rin106_32 in106_31 in106_32 9.241569
Rin106_33 in106_32 in106_33 9.241569
Rin106_34 in106_33 in106_34 9.241569
Rin106_35 in106_34 in106_35 9.241569
Rin106_36 in106_35 in106_36 9.241569
Rin106_37 in106_36 in106_37 9.241569
Rin106_38 in106_37 in106_38 9.241569
Rin106_39 in106_38 in106_39 9.241569
Rin106_40 in106_39 in106_40 9.241569
Rin106_41 in106_40 in106_41 9.241569
Rin106_42 in106_41 in106_42 9.241569
Rin106_43 in106_42 in106_43 9.241569
Rin106_44 in106_43 in106_44 9.241569
Rin106_45 in106_44 in106_45 9.241569
Rin106_46 in106_45 in106_46 9.241569
Rin106_47 in106_46 in106_47 9.241569
Rin106_48 in106_47 in106_48 9.241569
Rin106_49 in106_48 in106_49 9.241569
Rin106_50 in106_49 in106_50 9.241569
Rin106_51 in106_50 in106_51 9.241569
Rin106_52 in106_51 in106_52 9.241569
Rin106_53 in106_52 in106_53 9.241569
Rin106_54 in106_53 in106_54 9.241569
Rin106_55 in106_54 in106_55 9.241569
Rin106_56 in106_55 in106_56 9.241569
Rin106_57 in106 in106_57 9.241569
Rin106_58 in106_57 in106_58 9.241569
Rin106_59 in106_58 in106_59 9.241569
Rin106_60 in106_59 in106_60 9.241569
Rin106_61 in106_60 in106_61 9.241569
Rin106_62 in106_61 in106_62 9.241569
Rin106_63 in106_62 in106_63 9.241569
Rin106_64 in106_63 in106_64 9.241569
Rin106_65 in106_64 in106_65 9.241569
Rin106_66 in106_65 in106_66 9.241569
Rin106_67 in106_66 in106_67 9.241569
Rin106_68 in106_67 in106_68 9.241569
Rin106_69 in106_68 in106_69 9.241569
Rin106_70 in106_69 in106_70 9.241569
Rin106_71 in106_70 in106_71 9.241569
Rin106_72 in106_71 in106_72 9.241569
Rin106_73 in106_72 in106_73 9.241569
Rin106_74 in106_73 in106_74 9.241569
Rin106_75 in106_74 in106_75 9.241569
Rin106_76 in106_75 in106_76 9.241569
Rin106_77 in106_76 in106_77 9.241569
Rin106_78 in106_77 in106_78 9.241569
Rin106_79 in106_78 in106_79 9.241569
Rin106_80 in106_79 in106_80 9.241569
Rin106_81 in106_80 in106_81 9.241569
Rin106_82 in106_81 in106_82 9.241569
Rin106_83 in106_82 in106_83 9.241569
Rin106_84 in106_83 in106_84 9.241569
Rin107_1 in107 in107_1 9.241569
Rin107_2 in107_1 in107_2 9.241569
Rin107_3 in107_2 in107_3 9.241569
Rin107_4 in107_3 in107_4 9.241569
Rin107_5 in107_4 in107_5 9.241569
Rin107_6 in107_5 in107_6 9.241569
Rin107_7 in107_6 in107_7 9.241569
Rin107_8 in107_7 in107_8 9.241569
Rin107_9 in107_8 in107_9 9.241569
Rin107_10 in107_9 in107_10 9.241569
Rin107_11 in107_10 in107_11 9.241569
Rin107_12 in107_11 in107_12 9.241569
Rin107_13 in107_12 in107_13 9.241569
Rin107_14 in107_13 in107_14 9.241569
Rin107_15 in107_14 in107_15 9.241569
Rin107_16 in107_15 in107_16 9.241569
Rin107_17 in107_16 in107_17 9.241569
Rin107_18 in107_17 in107_18 9.241569
Rin107_19 in107_18 in107_19 9.241569
Rin107_20 in107_19 in107_20 9.241569
Rin107_21 in107_20 in107_21 9.241569
Rin107_22 in107_21 in107_22 9.241569
Rin107_23 in107_22 in107_23 9.241569
Rin107_24 in107_23 in107_24 9.241569
Rin107_25 in107_24 in107_25 9.241569
Rin107_26 in107_25 in107_26 9.241569
Rin107_27 in107_26 in107_27 9.241569
Rin107_28 in107_27 in107_28 9.241569
Rin107_29 in107 in107_29 9.241569
Rin107_30 in107_29 in107_30 9.241569
Rin107_31 in107_30 in107_31 9.241569
Rin107_32 in107_31 in107_32 9.241569
Rin107_33 in107_32 in107_33 9.241569
Rin107_34 in107_33 in107_34 9.241569
Rin107_35 in107_34 in107_35 9.241569
Rin107_36 in107_35 in107_36 9.241569
Rin107_37 in107_36 in107_37 9.241569
Rin107_38 in107_37 in107_38 9.241569
Rin107_39 in107_38 in107_39 9.241569
Rin107_40 in107_39 in107_40 9.241569
Rin107_41 in107_40 in107_41 9.241569
Rin107_42 in107_41 in107_42 9.241569
Rin107_43 in107_42 in107_43 9.241569
Rin107_44 in107_43 in107_44 9.241569
Rin107_45 in107_44 in107_45 9.241569
Rin107_46 in107_45 in107_46 9.241569
Rin107_47 in107_46 in107_47 9.241569
Rin107_48 in107_47 in107_48 9.241569
Rin107_49 in107_48 in107_49 9.241569
Rin107_50 in107_49 in107_50 9.241569
Rin107_51 in107_50 in107_51 9.241569
Rin107_52 in107_51 in107_52 9.241569
Rin107_53 in107_52 in107_53 9.241569
Rin107_54 in107_53 in107_54 9.241569
Rin107_55 in107_54 in107_55 9.241569
Rin107_56 in107_55 in107_56 9.241569
Rin107_57 in107 in107_57 9.241569
Rin107_58 in107_57 in107_58 9.241569
Rin107_59 in107_58 in107_59 9.241569
Rin107_60 in107_59 in107_60 9.241569
Rin107_61 in107_60 in107_61 9.241569
Rin107_62 in107_61 in107_62 9.241569
Rin107_63 in107_62 in107_63 9.241569
Rin107_64 in107_63 in107_64 9.241569
Rin107_65 in107_64 in107_65 9.241569
Rin107_66 in107_65 in107_66 9.241569
Rin107_67 in107_66 in107_67 9.241569
Rin107_68 in107_67 in107_68 9.241569
Rin107_69 in107_68 in107_69 9.241569
Rin107_70 in107_69 in107_70 9.241569
Rin107_71 in107_70 in107_71 9.241569
Rin107_72 in107_71 in107_72 9.241569
Rin107_73 in107_72 in107_73 9.241569
Rin107_74 in107_73 in107_74 9.241569
Rin107_75 in107_74 in107_75 9.241569
Rin107_76 in107_75 in107_76 9.241569
Rin107_77 in107_76 in107_77 9.241569
Rin107_78 in107_77 in107_78 9.241569
Rin107_79 in107_78 in107_79 9.241569
Rin107_80 in107_79 in107_80 9.241569
Rin107_81 in107_80 in107_81 9.241569
Rin107_82 in107_81 in107_82 9.241569
Rin107_83 in107_82 in107_83 9.241569
Rin107_84 in107_83 in107_84 9.241569
Rin108_1 in108 in108_1 9.241569
Rin108_2 in108_1 in108_2 9.241569
Rin108_3 in108_2 in108_3 9.241569
Rin108_4 in108_3 in108_4 9.241569
Rin108_5 in108_4 in108_5 9.241569
Rin108_6 in108_5 in108_6 9.241569
Rin108_7 in108_6 in108_7 9.241569
Rin108_8 in108_7 in108_8 9.241569
Rin108_9 in108_8 in108_9 9.241569
Rin108_10 in108_9 in108_10 9.241569
Rin108_11 in108_10 in108_11 9.241569
Rin108_12 in108_11 in108_12 9.241569
Rin108_13 in108_12 in108_13 9.241569
Rin108_14 in108_13 in108_14 9.241569
Rin108_15 in108_14 in108_15 9.241569
Rin108_16 in108_15 in108_16 9.241569
Rin108_17 in108_16 in108_17 9.241569
Rin108_18 in108_17 in108_18 9.241569
Rin108_19 in108_18 in108_19 9.241569
Rin108_20 in108_19 in108_20 9.241569
Rin108_21 in108_20 in108_21 9.241569
Rin108_22 in108_21 in108_22 9.241569
Rin108_23 in108_22 in108_23 9.241569
Rin108_24 in108_23 in108_24 9.241569
Rin108_25 in108_24 in108_25 9.241569
Rin108_26 in108_25 in108_26 9.241569
Rin108_27 in108_26 in108_27 9.241569
Rin108_28 in108_27 in108_28 9.241569
Rin108_29 in108 in108_29 9.241569
Rin108_30 in108_29 in108_30 9.241569
Rin108_31 in108_30 in108_31 9.241569
Rin108_32 in108_31 in108_32 9.241569
Rin108_33 in108_32 in108_33 9.241569
Rin108_34 in108_33 in108_34 9.241569
Rin108_35 in108_34 in108_35 9.241569
Rin108_36 in108_35 in108_36 9.241569
Rin108_37 in108_36 in108_37 9.241569
Rin108_38 in108_37 in108_38 9.241569
Rin108_39 in108_38 in108_39 9.241569
Rin108_40 in108_39 in108_40 9.241569
Rin108_41 in108_40 in108_41 9.241569
Rin108_42 in108_41 in108_42 9.241569
Rin108_43 in108_42 in108_43 9.241569
Rin108_44 in108_43 in108_44 9.241569
Rin108_45 in108_44 in108_45 9.241569
Rin108_46 in108_45 in108_46 9.241569
Rin108_47 in108_46 in108_47 9.241569
Rin108_48 in108_47 in108_48 9.241569
Rin108_49 in108_48 in108_49 9.241569
Rin108_50 in108_49 in108_50 9.241569
Rin108_51 in108_50 in108_51 9.241569
Rin108_52 in108_51 in108_52 9.241569
Rin108_53 in108_52 in108_53 9.241569
Rin108_54 in108_53 in108_54 9.241569
Rin108_55 in108_54 in108_55 9.241569
Rin108_56 in108_55 in108_56 9.241569
Rin108_57 in108 in108_57 9.241569
Rin108_58 in108_57 in108_58 9.241569
Rin108_59 in108_58 in108_59 9.241569
Rin108_60 in108_59 in108_60 9.241569
Rin108_61 in108_60 in108_61 9.241569
Rin108_62 in108_61 in108_62 9.241569
Rin108_63 in108_62 in108_63 9.241569
Rin108_64 in108_63 in108_64 9.241569
Rin108_65 in108_64 in108_65 9.241569
Rin108_66 in108_65 in108_66 9.241569
Rin108_67 in108_66 in108_67 9.241569
Rin108_68 in108_67 in108_68 9.241569
Rin108_69 in108_68 in108_69 9.241569
Rin108_70 in108_69 in108_70 9.241569
Rin108_71 in108_70 in108_71 9.241569
Rin108_72 in108_71 in108_72 9.241569
Rin108_73 in108_72 in108_73 9.241569
Rin108_74 in108_73 in108_74 9.241569
Rin108_75 in108_74 in108_75 9.241569
Rin108_76 in108_75 in108_76 9.241569
Rin108_77 in108_76 in108_77 9.241569
Rin108_78 in108_77 in108_78 9.241569
Rin108_79 in108_78 in108_79 9.241569
Rin108_80 in108_79 in108_80 9.241569
Rin108_81 in108_80 in108_81 9.241569
Rin108_82 in108_81 in108_82 9.241569
Rin108_83 in108_82 in108_83 9.241569
Rin108_84 in108_83 in108_84 9.241569
Rin109_1 in109 in109_1 9.241569
Rin109_2 in109_1 in109_2 9.241569
Rin109_3 in109_2 in109_3 9.241569
Rin109_4 in109_3 in109_4 9.241569
Rin109_5 in109_4 in109_5 9.241569
Rin109_6 in109_5 in109_6 9.241569
Rin109_7 in109_6 in109_7 9.241569
Rin109_8 in109_7 in109_8 9.241569
Rin109_9 in109_8 in109_9 9.241569
Rin109_10 in109_9 in109_10 9.241569
Rin109_11 in109_10 in109_11 9.241569
Rin109_12 in109_11 in109_12 9.241569
Rin109_13 in109_12 in109_13 9.241569
Rin109_14 in109_13 in109_14 9.241569
Rin109_15 in109_14 in109_15 9.241569
Rin109_16 in109_15 in109_16 9.241569
Rin109_17 in109_16 in109_17 9.241569
Rin109_18 in109_17 in109_18 9.241569
Rin109_19 in109_18 in109_19 9.241569
Rin109_20 in109_19 in109_20 9.241569
Rin109_21 in109_20 in109_21 9.241569
Rin109_22 in109_21 in109_22 9.241569
Rin109_23 in109_22 in109_23 9.241569
Rin109_24 in109_23 in109_24 9.241569
Rin109_25 in109_24 in109_25 9.241569
Rin109_26 in109_25 in109_26 9.241569
Rin109_27 in109_26 in109_27 9.241569
Rin109_28 in109_27 in109_28 9.241569
Rin109_29 in109 in109_29 9.241569
Rin109_30 in109_29 in109_30 9.241569
Rin109_31 in109_30 in109_31 9.241569
Rin109_32 in109_31 in109_32 9.241569
Rin109_33 in109_32 in109_33 9.241569
Rin109_34 in109_33 in109_34 9.241569
Rin109_35 in109_34 in109_35 9.241569
Rin109_36 in109_35 in109_36 9.241569
Rin109_37 in109_36 in109_37 9.241569
Rin109_38 in109_37 in109_38 9.241569
Rin109_39 in109_38 in109_39 9.241569
Rin109_40 in109_39 in109_40 9.241569
Rin109_41 in109_40 in109_41 9.241569
Rin109_42 in109_41 in109_42 9.241569
Rin109_43 in109_42 in109_43 9.241569
Rin109_44 in109_43 in109_44 9.241569
Rin109_45 in109_44 in109_45 9.241569
Rin109_46 in109_45 in109_46 9.241569
Rin109_47 in109_46 in109_47 9.241569
Rin109_48 in109_47 in109_48 9.241569
Rin109_49 in109_48 in109_49 9.241569
Rin109_50 in109_49 in109_50 9.241569
Rin109_51 in109_50 in109_51 9.241569
Rin109_52 in109_51 in109_52 9.241569
Rin109_53 in109_52 in109_53 9.241569
Rin109_54 in109_53 in109_54 9.241569
Rin109_55 in109_54 in109_55 9.241569
Rin109_56 in109_55 in109_56 9.241569
Rin109_57 in109 in109_57 9.241569
Rin109_58 in109_57 in109_58 9.241569
Rin109_59 in109_58 in109_59 9.241569
Rin109_60 in109_59 in109_60 9.241569
Rin109_61 in109_60 in109_61 9.241569
Rin109_62 in109_61 in109_62 9.241569
Rin109_63 in109_62 in109_63 9.241569
Rin109_64 in109_63 in109_64 9.241569
Rin109_65 in109_64 in109_65 9.241569
Rin109_66 in109_65 in109_66 9.241569
Rin109_67 in109_66 in109_67 9.241569
Rin109_68 in109_67 in109_68 9.241569
Rin109_69 in109_68 in109_69 9.241569
Rin109_70 in109_69 in109_70 9.241569
Rin109_71 in109_70 in109_71 9.241569
Rin109_72 in109_71 in109_72 9.241569
Rin109_73 in109_72 in109_73 9.241569
Rin109_74 in109_73 in109_74 9.241569
Rin109_75 in109_74 in109_75 9.241569
Rin109_76 in109_75 in109_76 9.241569
Rin109_77 in109_76 in109_77 9.241569
Rin109_78 in109_77 in109_78 9.241569
Rin109_79 in109_78 in109_79 9.241569
Rin109_80 in109_79 in109_80 9.241569
Rin109_81 in109_80 in109_81 9.241569
Rin109_82 in109_81 in109_82 9.241569
Rin109_83 in109_82 in109_83 9.241569
Rin109_84 in109_83 in109_84 9.241569
Rin110_1 in110 in110_1 9.241569
Rin110_2 in110_1 in110_2 9.241569
Rin110_3 in110_2 in110_3 9.241569
Rin110_4 in110_3 in110_4 9.241569
Rin110_5 in110_4 in110_5 9.241569
Rin110_6 in110_5 in110_6 9.241569
Rin110_7 in110_6 in110_7 9.241569
Rin110_8 in110_7 in110_8 9.241569
Rin110_9 in110_8 in110_9 9.241569
Rin110_10 in110_9 in110_10 9.241569
Rin110_11 in110_10 in110_11 9.241569
Rin110_12 in110_11 in110_12 9.241569
Rin110_13 in110_12 in110_13 9.241569
Rin110_14 in110_13 in110_14 9.241569
Rin110_15 in110_14 in110_15 9.241569
Rin110_16 in110_15 in110_16 9.241569
Rin110_17 in110_16 in110_17 9.241569
Rin110_18 in110_17 in110_18 9.241569
Rin110_19 in110_18 in110_19 9.241569
Rin110_20 in110_19 in110_20 9.241569
Rin110_21 in110_20 in110_21 9.241569
Rin110_22 in110_21 in110_22 9.241569
Rin110_23 in110_22 in110_23 9.241569
Rin110_24 in110_23 in110_24 9.241569
Rin110_25 in110_24 in110_25 9.241569
Rin110_26 in110_25 in110_26 9.241569
Rin110_27 in110_26 in110_27 9.241569
Rin110_28 in110_27 in110_28 9.241569
Rin110_29 in110 in110_29 9.241569
Rin110_30 in110_29 in110_30 9.241569
Rin110_31 in110_30 in110_31 9.241569
Rin110_32 in110_31 in110_32 9.241569
Rin110_33 in110_32 in110_33 9.241569
Rin110_34 in110_33 in110_34 9.241569
Rin110_35 in110_34 in110_35 9.241569
Rin110_36 in110_35 in110_36 9.241569
Rin110_37 in110_36 in110_37 9.241569
Rin110_38 in110_37 in110_38 9.241569
Rin110_39 in110_38 in110_39 9.241569
Rin110_40 in110_39 in110_40 9.241569
Rin110_41 in110_40 in110_41 9.241569
Rin110_42 in110_41 in110_42 9.241569
Rin110_43 in110_42 in110_43 9.241569
Rin110_44 in110_43 in110_44 9.241569
Rin110_45 in110_44 in110_45 9.241569
Rin110_46 in110_45 in110_46 9.241569
Rin110_47 in110_46 in110_47 9.241569
Rin110_48 in110_47 in110_48 9.241569
Rin110_49 in110_48 in110_49 9.241569
Rin110_50 in110_49 in110_50 9.241569
Rin110_51 in110_50 in110_51 9.241569
Rin110_52 in110_51 in110_52 9.241569
Rin110_53 in110_52 in110_53 9.241569
Rin110_54 in110_53 in110_54 9.241569
Rin110_55 in110_54 in110_55 9.241569
Rin110_56 in110_55 in110_56 9.241569
Rin110_57 in110 in110_57 9.241569
Rin110_58 in110_57 in110_58 9.241569
Rin110_59 in110_58 in110_59 9.241569
Rin110_60 in110_59 in110_60 9.241569
Rin110_61 in110_60 in110_61 9.241569
Rin110_62 in110_61 in110_62 9.241569
Rin110_63 in110_62 in110_63 9.241569
Rin110_64 in110_63 in110_64 9.241569
Rin110_65 in110_64 in110_65 9.241569
Rin110_66 in110_65 in110_66 9.241569
Rin110_67 in110_66 in110_67 9.241569
Rin110_68 in110_67 in110_68 9.241569
Rin110_69 in110_68 in110_69 9.241569
Rin110_70 in110_69 in110_70 9.241569
Rin110_71 in110_70 in110_71 9.241569
Rin110_72 in110_71 in110_72 9.241569
Rin110_73 in110_72 in110_73 9.241569
Rin110_74 in110_73 in110_74 9.241569
Rin110_75 in110_74 in110_75 9.241569
Rin110_76 in110_75 in110_76 9.241569
Rin110_77 in110_76 in110_77 9.241569
Rin110_78 in110_77 in110_78 9.241569
Rin110_79 in110_78 in110_79 9.241569
Rin110_80 in110_79 in110_80 9.241569
Rin110_81 in110_80 in110_81 9.241569
Rin110_82 in110_81 in110_82 9.241569
Rin110_83 in110_82 in110_83 9.241569
Rin110_84 in110_83 in110_84 9.241569
Rin111_1 in111 in111_1 9.241569
Rin111_2 in111_1 in111_2 9.241569
Rin111_3 in111_2 in111_3 9.241569
Rin111_4 in111_3 in111_4 9.241569
Rin111_5 in111_4 in111_5 9.241569
Rin111_6 in111_5 in111_6 9.241569
Rin111_7 in111_6 in111_7 9.241569
Rin111_8 in111_7 in111_8 9.241569
Rin111_9 in111_8 in111_9 9.241569
Rin111_10 in111_9 in111_10 9.241569
Rin111_11 in111_10 in111_11 9.241569
Rin111_12 in111_11 in111_12 9.241569
Rin111_13 in111_12 in111_13 9.241569
Rin111_14 in111_13 in111_14 9.241569
Rin111_15 in111_14 in111_15 9.241569
Rin111_16 in111_15 in111_16 9.241569
Rin111_17 in111_16 in111_17 9.241569
Rin111_18 in111_17 in111_18 9.241569
Rin111_19 in111_18 in111_19 9.241569
Rin111_20 in111_19 in111_20 9.241569
Rin111_21 in111_20 in111_21 9.241569
Rin111_22 in111_21 in111_22 9.241569
Rin111_23 in111_22 in111_23 9.241569
Rin111_24 in111_23 in111_24 9.241569
Rin111_25 in111_24 in111_25 9.241569
Rin111_26 in111_25 in111_26 9.241569
Rin111_27 in111_26 in111_27 9.241569
Rin111_28 in111_27 in111_28 9.241569
Rin111_29 in111 in111_29 9.241569
Rin111_30 in111_29 in111_30 9.241569
Rin111_31 in111_30 in111_31 9.241569
Rin111_32 in111_31 in111_32 9.241569
Rin111_33 in111_32 in111_33 9.241569
Rin111_34 in111_33 in111_34 9.241569
Rin111_35 in111_34 in111_35 9.241569
Rin111_36 in111_35 in111_36 9.241569
Rin111_37 in111_36 in111_37 9.241569
Rin111_38 in111_37 in111_38 9.241569
Rin111_39 in111_38 in111_39 9.241569
Rin111_40 in111_39 in111_40 9.241569
Rin111_41 in111_40 in111_41 9.241569
Rin111_42 in111_41 in111_42 9.241569
Rin111_43 in111_42 in111_43 9.241569
Rin111_44 in111_43 in111_44 9.241569
Rin111_45 in111_44 in111_45 9.241569
Rin111_46 in111_45 in111_46 9.241569
Rin111_47 in111_46 in111_47 9.241569
Rin111_48 in111_47 in111_48 9.241569
Rin111_49 in111_48 in111_49 9.241569
Rin111_50 in111_49 in111_50 9.241569
Rin111_51 in111_50 in111_51 9.241569
Rin111_52 in111_51 in111_52 9.241569
Rin111_53 in111_52 in111_53 9.241569
Rin111_54 in111_53 in111_54 9.241569
Rin111_55 in111_54 in111_55 9.241569
Rin111_56 in111_55 in111_56 9.241569
Rin111_57 in111 in111_57 9.241569
Rin111_58 in111_57 in111_58 9.241569
Rin111_59 in111_58 in111_59 9.241569
Rin111_60 in111_59 in111_60 9.241569
Rin111_61 in111_60 in111_61 9.241569
Rin111_62 in111_61 in111_62 9.241569
Rin111_63 in111_62 in111_63 9.241569
Rin111_64 in111_63 in111_64 9.241569
Rin111_65 in111_64 in111_65 9.241569
Rin111_66 in111_65 in111_66 9.241569
Rin111_67 in111_66 in111_67 9.241569
Rin111_68 in111_67 in111_68 9.241569
Rin111_69 in111_68 in111_69 9.241569
Rin111_70 in111_69 in111_70 9.241569
Rin111_71 in111_70 in111_71 9.241569
Rin111_72 in111_71 in111_72 9.241569
Rin111_73 in111_72 in111_73 9.241569
Rin111_74 in111_73 in111_74 9.241569
Rin111_75 in111_74 in111_75 9.241569
Rin111_76 in111_75 in111_76 9.241569
Rin111_77 in111_76 in111_77 9.241569
Rin111_78 in111_77 in111_78 9.241569
Rin111_79 in111_78 in111_79 9.241569
Rin111_80 in111_79 in111_80 9.241569
Rin111_81 in111_80 in111_81 9.241569
Rin111_82 in111_81 in111_82 9.241569
Rin111_83 in111_82 in111_83 9.241569
Rin111_84 in111_83 in111_84 9.241569
Rin112_1 in112 in112_1 9.241569
Rin112_2 in112_1 in112_2 9.241569
Rin112_3 in112_2 in112_3 9.241569
Rin112_4 in112_3 in112_4 9.241569
Rin112_5 in112_4 in112_5 9.241569
Rin112_6 in112_5 in112_6 9.241569
Rin112_7 in112_6 in112_7 9.241569
Rin112_8 in112_7 in112_8 9.241569
Rin112_9 in112_8 in112_9 9.241569
Rin112_10 in112_9 in112_10 9.241569
Rin112_11 in112_10 in112_11 9.241569
Rin112_12 in112_11 in112_12 9.241569
Rin112_13 in112_12 in112_13 9.241569
Rin112_14 in112_13 in112_14 9.241569
Rin112_15 in112_14 in112_15 9.241569
Rin112_16 in112_15 in112_16 9.241569
Rin112_17 in112_16 in112_17 9.241569
Rin112_18 in112_17 in112_18 9.241569
Rin112_19 in112_18 in112_19 9.241569
Rin112_20 in112_19 in112_20 9.241569
Rin112_21 in112_20 in112_21 9.241569
Rin112_22 in112_21 in112_22 9.241569
Rin112_23 in112_22 in112_23 9.241569
Rin112_24 in112_23 in112_24 9.241569
Rin112_25 in112_24 in112_25 9.241569
Rin112_26 in112_25 in112_26 9.241569
Rin112_27 in112_26 in112_27 9.241569
Rin112_28 in112_27 in112_28 9.241569
Rin112_29 in112 in112_29 9.241569
Rin112_30 in112_29 in112_30 9.241569
Rin112_31 in112_30 in112_31 9.241569
Rin112_32 in112_31 in112_32 9.241569
Rin112_33 in112_32 in112_33 9.241569
Rin112_34 in112_33 in112_34 9.241569
Rin112_35 in112_34 in112_35 9.241569
Rin112_36 in112_35 in112_36 9.241569
Rin112_37 in112_36 in112_37 9.241569
Rin112_38 in112_37 in112_38 9.241569
Rin112_39 in112_38 in112_39 9.241569
Rin112_40 in112_39 in112_40 9.241569
Rin112_41 in112_40 in112_41 9.241569
Rin112_42 in112_41 in112_42 9.241569
Rin112_43 in112_42 in112_43 9.241569
Rin112_44 in112_43 in112_44 9.241569
Rin112_45 in112_44 in112_45 9.241569
Rin112_46 in112_45 in112_46 9.241569
Rin112_47 in112_46 in112_47 9.241569
Rin112_48 in112_47 in112_48 9.241569
Rin112_49 in112_48 in112_49 9.241569
Rin112_50 in112_49 in112_50 9.241569
Rin112_51 in112_50 in112_51 9.241569
Rin112_52 in112_51 in112_52 9.241569
Rin112_53 in112_52 in112_53 9.241569
Rin112_54 in112_53 in112_54 9.241569
Rin112_55 in112_54 in112_55 9.241569
Rin112_56 in112_55 in112_56 9.241569
Rin112_57 in112 in112_57 9.241569
Rin112_58 in112_57 in112_58 9.241569
Rin112_59 in112_58 in112_59 9.241569
Rin112_60 in112_59 in112_60 9.241569
Rin112_61 in112_60 in112_61 9.241569
Rin112_62 in112_61 in112_62 9.241569
Rin112_63 in112_62 in112_63 9.241569
Rin112_64 in112_63 in112_64 9.241569
Rin112_65 in112_64 in112_65 9.241569
Rin112_66 in112_65 in112_66 9.241569
Rin112_67 in112_66 in112_67 9.241569
Rin112_68 in112_67 in112_68 9.241569
Rin112_69 in112_68 in112_69 9.241569
Rin112_70 in112_69 in112_70 9.241569
Rin112_71 in112_70 in112_71 9.241569
Rin112_72 in112_71 in112_72 9.241569
Rin112_73 in112_72 in112_73 9.241569
Rin112_74 in112_73 in112_74 9.241569
Rin112_75 in112_74 in112_75 9.241569
Rin112_76 in112_75 in112_76 9.241569
Rin112_77 in112_76 in112_77 9.241569
Rin112_78 in112_77 in112_78 9.241569
Rin112_79 in112_78 in112_79 9.241569
Rin112_80 in112_79 in112_80 9.241569
Rin112_81 in112_80 in112_81 9.241569
Rin112_82 in112_81 in112_82 9.241569
Rin112_83 in112_82 in112_83 9.241569
Rin112_84 in112_83 in112_84 9.241569
Rin113_1 in113 in113_1 9.241569
Rin113_2 in113_1 in113_2 9.241569
Rin113_3 in113_2 in113_3 9.241569
Rin113_4 in113_3 in113_4 9.241569
Rin113_5 in113_4 in113_5 9.241569
Rin113_6 in113_5 in113_6 9.241569
Rin113_7 in113_6 in113_7 9.241569
Rin113_8 in113_7 in113_8 9.241569
Rin113_9 in113_8 in113_9 9.241569
Rin113_10 in113_9 in113_10 9.241569
Rin113_11 in113_10 in113_11 9.241569
Rin113_12 in113_11 in113_12 9.241569
Rin113_13 in113_12 in113_13 9.241569
Rin113_14 in113_13 in113_14 9.241569
Rin113_15 in113_14 in113_15 9.241569
Rin113_16 in113_15 in113_16 9.241569
Rin113_17 in113_16 in113_17 9.241569
Rin113_18 in113_17 in113_18 9.241569
Rin113_19 in113_18 in113_19 9.241569
Rin113_20 in113_19 in113_20 9.241569
Rin113_21 in113_20 in113_21 9.241569
Rin113_22 in113_21 in113_22 9.241569
Rin113_23 in113_22 in113_23 9.241569
Rin113_24 in113_23 in113_24 9.241569
Rin113_25 in113_24 in113_25 9.241569
Rin113_26 in113_25 in113_26 9.241569
Rin113_27 in113_26 in113_27 9.241569
Rin113_28 in113_27 in113_28 9.241569
Rin113_29 in113 in113_29 9.241569
Rin113_30 in113_29 in113_30 9.241569
Rin113_31 in113_30 in113_31 9.241569
Rin113_32 in113_31 in113_32 9.241569
Rin113_33 in113_32 in113_33 9.241569
Rin113_34 in113_33 in113_34 9.241569
Rin113_35 in113_34 in113_35 9.241569
Rin113_36 in113_35 in113_36 9.241569
Rin113_37 in113_36 in113_37 9.241569
Rin113_38 in113_37 in113_38 9.241569
Rin113_39 in113_38 in113_39 9.241569
Rin113_40 in113_39 in113_40 9.241569
Rin113_41 in113_40 in113_41 9.241569
Rin113_42 in113_41 in113_42 9.241569
Rin113_43 in113_42 in113_43 9.241569
Rin113_44 in113_43 in113_44 9.241569
Rin113_45 in113_44 in113_45 9.241569
Rin113_46 in113_45 in113_46 9.241569
Rin113_47 in113_46 in113_47 9.241569
Rin113_48 in113_47 in113_48 9.241569
Rin113_49 in113_48 in113_49 9.241569
Rin113_50 in113_49 in113_50 9.241569
Rin113_51 in113_50 in113_51 9.241569
Rin113_52 in113_51 in113_52 9.241569
Rin113_53 in113_52 in113_53 9.241569
Rin113_54 in113_53 in113_54 9.241569
Rin113_55 in113_54 in113_55 9.241569
Rin113_56 in113_55 in113_56 9.241569
Rin113_57 in113 in113_57 9.241569
Rin113_58 in113_57 in113_58 9.241569
Rin113_59 in113_58 in113_59 9.241569
Rin113_60 in113_59 in113_60 9.241569
Rin113_61 in113_60 in113_61 9.241569
Rin113_62 in113_61 in113_62 9.241569
Rin113_63 in113_62 in113_63 9.241569
Rin113_64 in113_63 in113_64 9.241569
Rin113_65 in113_64 in113_65 9.241569
Rin113_66 in113_65 in113_66 9.241569
Rin113_67 in113_66 in113_67 9.241569
Rin113_68 in113_67 in113_68 9.241569
Rin113_69 in113_68 in113_69 9.241569
Rin113_70 in113_69 in113_70 9.241569
Rin113_71 in113_70 in113_71 9.241569
Rin113_72 in113_71 in113_72 9.241569
Rin113_73 in113_72 in113_73 9.241569
Rin113_74 in113_73 in113_74 9.241569
Rin113_75 in113_74 in113_75 9.241569
Rin113_76 in113_75 in113_76 9.241569
Rin113_77 in113_76 in113_77 9.241569
Rin113_78 in113_77 in113_78 9.241569
Rin113_79 in113_78 in113_79 9.241569
Rin113_80 in113_79 in113_80 9.241569
Rin113_81 in113_80 in113_81 9.241569
Rin113_82 in113_81 in113_82 9.241569
Rin113_83 in113_82 in113_83 9.241569
Rin113_84 in113_83 in113_84 9.241569
Rin114_1 in114 in114_1 9.241569
Rin114_2 in114_1 in114_2 9.241569
Rin114_3 in114_2 in114_3 9.241569
Rin114_4 in114_3 in114_4 9.241569
Rin114_5 in114_4 in114_5 9.241569
Rin114_6 in114_5 in114_6 9.241569
Rin114_7 in114_6 in114_7 9.241569
Rin114_8 in114_7 in114_8 9.241569
Rin114_9 in114_8 in114_9 9.241569
Rin114_10 in114_9 in114_10 9.241569
Rin114_11 in114_10 in114_11 9.241569
Rin114_12 in114_11 in114_12 9.241569
Rin114_13 in114_12 in114_13 9.241569
Rin114_14 in114_13 in114_14 9.241569
Rin114_15 in114_14 in114_15 9.241569
Rin114_16 in114_15 in114_16 9.241569
Rin114_17 in114_16 in114_17 9.241569
Rin114_18 in114_17 in114_18 9.241569
Rin114_19 in114_18 in114_19 9.241569
Rin114_20 in114_19 in114_20 9.241569
Rin114_21 in114_20 in114_21 9.241569
Rin114_22 in114_21 in114_22 9.241569
Rin114_23 in114_22 in114_23 9.241569
Rin114_24 in114_23 in114_24 9.241569
Rin114_25 in114_24 in114_25 9.241569
Rin114_26 in114_25 in114_26 9.241569
Rin114_27 in114_26 in114_27 9.241569
Rin114_28 in114_27 in114_28 9.241569
Rin114_29 in114 in114_29 9.241569
Rin114_30 in114_29 in114_30 9.241569
Rin114_31 in114_30 in114_31 9.241569
Rin114_32 in114_31 in114_32 9.241569
Rin114_33 in114_32 in114_33 9.241569
Rin114_34 in114_33 in114_34 9.241569
Rin114_35 in114_34 in114_35 9.241569
Rin114_36 in114_35 in114_36 9.241569
Rin114_37 in114_36 in114_37 9.241569
Rin114_38 in114_37 in114_38 9.241569
Rin114_39 in114_38 in114_39 9.241569
Rin114_40 in114_39 in114_40 9.241569
Rin114_41 in114_40 in114_41 9.241569
Rin114_42 in114_41 in114_42 9.241569
Rin114_43 in114_42 in114_43 9.241569
Rin114_44 in114_43 in114_44 9.241569
Rin114_45 in114_44 in114_45 9.241569
Rin114_46 in114_45 in114_46 9.241569
Rin114_47 in114_46 in114_47 9.241569
Rin114_48 in114_47 in114_48 9.241569
Rin114_49 in114_48 in114_49 9.241569
Rin114_50 in114_49 in114_50 9.241569
Rin114_51 in114_50 in114_51 9.241569
Rin114_52 in114_51 in114_52 9.241569
Rin114_53 in114_52 in114_53 9.241569
Rin114_54 in114_53 in114_54 9.241569
Rin114_55 in114_54 in114_55 9.241569
Rin114_56 in114_55 in114_56 9.241569
Rin114_57 in114 in114_57 9.241569
Rin114_58 in114_57 in114_58 9.241569
Rin114_59 in114_58 in114_59 9.241569
Rin114_60 in114_59 in114_60 9.241569
Rin114_61 in114_60 in114_61 9.241569
Rin114_62 in114_61 in114_62 9.241569
Rin114_63 in114_62 in114_63 9.241569
Rin114_64 in114_63 in114_64 9.241569
Rin114_65 in114_64 in114_65 9.241569
Rin114_66 in114_65 in114_66 9.241569
Rin114_67 in114_66 in114_67 9.241569
Rin114_68 in114_67 in114_68 9.241569
Rin114_69 in114_68 in114_69 9.241569
Rin114_70 in114_69 in114_70 9.241569
Rin114_71 in114_70 in114_71 9.241569
Rin114_72 in114_71 in114_72 9.241569
Rin114_73 in114_72 in114_73 9.241569
Rin114_74 in114_73 in114_74 9.241569
Rin114_75 in114_74 in114_75 9.241569
Rin114_76 in114_75 in114_76 9.241569
Rin114_77 in114_76 in114_77 9.241569
Rin114_78 in114_77 in114_78 9.241569
Rin114_79 in114_78 in114_79 9.241569
Rin114_80 in114_79 in114_80 9.241569
Rin114_81 in114_80 in114_81 9.241569
Rin114_82 in114_81 in114_82 9.241569
Rin114_83 in114_82 in114_83 9.241569
Rin114_84 in114_83 in114_84 9.241569
Rin115_1 in115 in115_1 9.241569
Rin115_2 in115_1 in115_2 9.241569
Rin115_3 in115_2 in115_3 9.241569
Rin115_4 in115_3 in115_4 9.241569
Rin115_5 in115_4 in115_5 9.241569
Rin115_6 in115_5 in115_6 9.241569
Rin115_7 in115_6 in115_7 9.241569
Rin115_8 in115_7 in115_8 9.241569
Rin115_9 in115_8 in115_9 9.241569
Rin115_10 in115_9 in115_10 9.241569
Rin115_11 in115_10 in115_11 9.241569
Rin115_12 in115_11 in115_12 9.241569
Rin115_13 in115_12 in115_13 9.241569
Rin115_14 in115_13 in115_14 9.241569
Rin115_15 in115_14 in115_15 9.241569
Rin115_16 in115_15 in115_16 9.241569
Rin115_17 in115_16 in115_17 9.241569
Rin115_18 in115_17 in115_18 9.241569
Rin115_19 in115_18 in115_19 9.241569
Rin115_20 in115_19 in115_20 9.241569
Rin115_21 in115_20 in115_21 9.241569
Rin115_22 in115_21 in115_22 9.241569
Rin115_23 in115_22 in115_23 9.241569
Rin115_24 in115_23 in115_24 9.241569
Rin115_25 in115_24 in115_25 9.241569
Rin115_26 in115_25 in115_26 9.241569
Rin115_27 in115_26 in115_27 9.241569
Rin115_28 in115_27 in115_28 9.241569
Rin115_29 in115 in115_29 9.241569
Rin115_30 in115_29 in115_30 9.241569
Rin115_31 in115_30 in115_31 9.241569
Rin115_32 in115_31 in115_32 9.241569
Rin115_33 in115_32 in115_33 9.241569
Rin115_34 in115_33 in115_34 9.241569
Rin115_35 in115_34 in115_35 9.241569
Rin115_36 in115_35 in115_36 9.241569
Rin115_37 in115_36 in115_37 9.241569
Rin115_38 in115_37 in115_38 9.241569
Rin115_39 in115_38 in115_39 9.241569
Rin115_40 in115_39 in115_40 9.241569
Rin115_41 in115_40 in115_41 9.241569
Rin115_42 in115_41 in115_42 9.241569
Rin115_43 in115_42 in115_43 9.241569
Rin115_44 in115_43 in115_44 9.241569
Rin115_45 in115_44 in115_45 9.241569
Rin115_46 in115_45 in115_46 9.241569
Rin115_47 in115_46 in115_47 9.241569
Rin115_48 in115_47 in115_48 9.241569
Rin115_49 in115_48 in115_49 9.241569
Rin115_50 in115_49 in115_50 9.241569
Rin115_51 in115_50 in115_51 9.241569
Rin115_52 in115_51 in115_52 9.241569
Rin115_53 in115_52 in115_53 9.241569
Rin115_54 in115_53 in115_54 9.241569
Rin115_55 in115_54 in115_55 9.241569
Rin115_56 in115_55 in115_56 9.241569
Rin115_57 in115 in115_57 9.241569
Rin115_58 in115_57 in115_58 9.241569
Rin115_59 in115_58 in115_59 9.241569
Rin115_60 in115_59 in115_60 9.241569
Rin115_61 in115_60 in115_61 9.241569
Rin115_62 in115_61 in115_62 9.241569
Rin115_63 in115_62 in115_63 9.241569
Rin115_64 in115_63 in115_64 9.241569
Rin115_65 in115_64 in115_65 9.241569
Rin115_66 in115_65 in115_66 9.241569
Rin115_67 in115_66 in115_67 9.241569
Rin115_68 in115_67 in115_68 9.241569
Rin115_69 in115_68 in115_69 9.241569
Rin115_70 in115_69 in115_70 9.241569
Rin115_71 in115_70 in115_71 9.241569
Rin115_72 in115_71 in115_72 9.241569
Rin115_73 in115_72 in115_73 9.241569
Rin115_74 in115_73 in115_74 9.241569
Rin115_75 in115_74 in115_75 9.241569
Rin115_76 in115_75 in115_76 9.241569
Rin115_77 in115_76 in115_77 9.241569
Rin115_78 in115_77 in115_78 9.241569
Rin115_79 in115_78 in115_79 9.241569
Rin115_80 in115_79 in115_80 9.241569
Rin115_81 in115_80 in115_81 9.241569
Rin115_82 in115_81 in115_82 9.241569
Rin115_83 in115_82 in115_83 9.241569
Rin115_84 in115_83 in115_84 9.241569
Rin116_1 in116 in116_1 9.241569
Rin116_2 in116_1 in116_2 9.241569
Rin116_3 in116_2 in116_3 9.241569
Rin116_4 in116_3 in116_4 9.241569
Rin116_5 in116_4 in116_5 9.241569
Rin116_6 in116_5 in116_6 9.241569
Rin116_7 in116_6 in116_7 9.241569
Rin116_8 in116_7 in116_8 9.241569
Rin116_9 in116_8 in116_9 9.241569
Rin116_10 in116_9 in116_10 9.241569
Rin116_11 in116_10 in116_11 9.241569
Rin116_12 in116_11 in116_12 9.241569
Rin116_13 in116_12 in116_13 9.241569
Rin116_14 in116_13 in116_14 9.241569
Rin116_15 in116_14 in116_15 9.241569
Rin116_16 in116_15 in116_16 9.241569
Rin116_17 in116_16 in116_17 9.241569
Rin116_18 in116_17 in116_18 9.241569
Rin116_19 in116_18 in116_19 9.241569
Rin116_20 in116_19 in116_20 9.241569
Rin116_21 in116_20 in116_21 9.241569
Rin116_22 in116_21 in116_22 9.241569
Rin116_23 in116_22 in116_23 9.241569
Rin116_24 in116_23 in116_24 9.241569
Rin116_25 in116_24 in116_25 9.241569
Rin116_26 in116_25 in116_26 9.241569
Rin116_27 in116_26 in116_27 9.241569
Rin116_28 in116_27 in116_28 9.241569
Rin116_29 in116 in116_29 9.241569
Rin116_30 in116_29 in116_30 9.241569
Rin116_31 in116_30 in116_31 9.241569
Rin116_32 in116_31 in116_32 9.241569
Rin116_33 in116_32 in116_33 9.241569
Rin116_34 in116_33 in116_34 9.241569
Rin116_35 in116_34 in116_35 9.241569
Rin116_36 in116_35 in116_36 9.241569
Rin116_37 in116_36 in116_37 9.241569
Rin116_38 in116_37 in116_38 9.241569
Rin116_39 in116_38 in116_39 9.241569
Rin116_40 in116_39 in116_40 9.241569
Rin116_41 in116_40 in116_41 9.241569
Rin116_42 in116_41 in116_42 9.241569
Rin116_43 in116_42 in116_43 9.241569
Rin116_44 in116_43 in116_44 9.241569
Rin116_45 in116_44 in116_45 9.241569
Rin116_46 in116_45 in116_46 9.241569
Rin116_47 in116_46 in116_47 9.241569
Rin116_48 in116_47 in116_48 9.241569
Rin116_49 in116_48 in116_49 9.241569
Rin116_50 in116_49 in116_50 9.241569
Rin116_51 in116_50 in116_51 9.241569
Rin116_52 in116_51 in116_52 9.241569
Rin116_53 in116_52 in116_53 9.241569
Rin116_54 in116_53 in116_54 9.241569
Rin116_55 in116_54 in116_55 9.241569
Rin116_56 in116_55 in116_56 9.241569
Rin116_57 in116 in116_57 9.241569
Rin116_58 in116_57 in116_58 9.241569
Rin116_59 in116_58 in116_59 9.241569
Rin116_60 in116_59 in116_60 9.241569
Rin116_61 in116_60 in116_61 9.241569
Rin116_62 in116_61 in116_62 9.241569
Rin116_63 in116_62 in116_63 9.241569
Rin116_64 in116_63 in116_64 9.241569
Rin116_65 in116_64 in116_65 9.241569
Rin116_66 in116_65 in116_66 9.241569
Rin116_67 in116_66 in116_67 9.241569
Rin116_68 in116_67 in116_68 9.241569
Rin116_69 in116_68 in116_69 9.241569
Rin116_70 in116_69 in116_70 9.241569
Rin116_71 in116_70 in116_71 9.241569
Rin116_72 in116_71 in116_72 9.241569
Rin116_73 in116_72 in116_73 9.241569
Rin116_74 in116_73 in116_74 9.241569
Rin116_75 in116_74 in116_75 9.241569
Rin116_76 in116_75 in116_76 9.241569
Rin116_77 in116_76 in116_77 9.241569
Rin116_78 in116_77 in116_78 9.241569
Rin116_79 in116_78 in116_79 9.241569
Rin116_80 in116_79 in116_80 9.241569
Rin116_81 in116_80 in116_81 9.241569
Rin116_82 in116_81 in116_82 9.241569
Rin116_83 in116_82 in116_83 9.241569
Rin116_84 in116_83 in116_84 9.241569
Rin117_1 in117 in117_1 9.241569
Rin117_2 in117_1 in117_2 9.241569
Rin117_3 in117_2 in117_3 9.241569
Rin117_4 in117_3 in117_4 9.241569
Rin117_5 in117_4 in117_5 9.241569
Rin117_6 in117_5 in117_6 9.241569
Rin117_7 in117_6 in117_7 9.241569
Rin117_8 in117_7 in117_8 9.241569
Rin117_9 in117_8 in117_9 9.241569
Rin117_10 in117_9 in117_10 9.241569
Rin117_11 in117_10 in117_11 9.241569
Rin117_12 in117_11 in117_12 9.241569
Rin117_13 in117_12 in117_13 9.241569
Rin117_14 in117_13 in117_14 9.241569
Rin117_15 in117_14 in117_15 9.241569
Rin117_16 in117_15 in117_16 9.241569
Rin117_17 in117_16 in117_17 9.241569
Rin117_18 in117_17 in117_18 9.241569
Rin117_19 in117_18 in117_19 9.241569
Rin117_20 in117_19 in117_20 9.241569
Rin117_21 in117_20 in117_21 9.241569
Rin117_22 in117_21 in117_22 9.241569
Rin117_23 in117_22 in117_23 9.241569
Rin117_24 in117_23 in117_24 9.241569
Rin117_25 in117_24 in117_25 9.241569
Rin117_26 in117_25 in117_26 9.241569
Rin117_27 in117_26 in117_27 9.241569
Rin117_28 in117_27 in117_28 9.241569
Rin117_29 in117 in117_29 9.241569
Rin117_30 in117_29 in117_30 9.241569
Rin117_31 in117_30 in117_31 9.241569
Rin117_32 in117_31 in117_32 9.241569
Rin117_33 in117_32 in117_33 9.241569
Rin117_34 in117_33 in117_34 9.241569
Rin117_35 in117_34 in117_35 9.241569
Rin117_36 in117_35 in117_36 9.241569
Rin117_37 in117_36 in117_37 9.241569
Rin117_38 in117_37 in117_38 9.241569
Rin117_39 in117_38 in117_39 9.241569
Rin117_40 in117_39 in117_40 9.241569
Rin117_41 in117_40 in117_41 9.241569
Rin117_42 in117_41 in117_42 9.241569
Rin117_43 in117_42 in117_43 9.241569
Rin117_44 in117_43 in117_44 9.241569
Rin117_45 in117_44 in117_45 9.241569
Rin117_46 in117_45 in117_46 9.241569
Rin117_47 in117_46 in117_47 9.241569
Rin117_48 in117_47 in117_48 9.241569
Rin117_49 in117_48 in117_49 9.241569
Rin117_50 in117_49 in117_50 9.241569
Rin117_51 in117_50 in117_51 9.241569
Rin117_52 in117_51 in117_52 9.241569
Rin117_53 in117_52 in117_53 9.241569
Rin117_54 in117_53 in117_54 9.241569
Rin117_55 in117_54 in117_55 9.241569
Rin117_56 in117_55 in117_56 9.241569
Rin117_57 in117 in117_57 9.241569
Rin117_58 in117_57 in117_58 9.241569
Rin117_59 in117_58 in117_59 9.241569
Rin117_60 in117_59 in117_60 9.241569
Rin117_61 in117_60 in117_61 9.241569
Rin117_62 in117_61 in117_62 9.241569
Rin117_63 in117_62 in117_63 9.241569
Rin117_64 in117_63 in117_64 9.241569
Rin117_65 in117_64 in117_65 9.241569
Rin117_66 in117_65 in117_66 9.241569
Rin117_67 in117_66 in117_67 9.241569
Rin117_68 in117_67 in117_68 9.241569
Rin117_69 in117_68 in117_69 9.241569
Rin117_70 in117_69 in117_70 9.241569
Rin117_71 in117_70 in117_71 9.241569
Rin117_72 in117_71 in117_72 9.241569
Rin117_73 in117_72 in117_73 9.241569
Rin117_74 in117_73 in117_74 9.241569
Rin117_75 in117_74 in117_75 9.241569
Rin117_76 in117_75 in117_76 9.241569
Rin117_77 in117_76 in117_77 9.241569
Rin117_78 in117_77 in117_78 9.241569
Rin117_79 in117_78 in117_79 9.241569
Rin117_80 in117_79 in117_80 9.241569
Rin117_81 in117_80 in117_81 9.241569
Rin117_82 in117_81 in117_82 9.241569
Rin117_83 in117_82 in117_83 9.241569
Rin117_84 in117_83 in117_84 9.241569
Rin118_1 in118 in118_1 9.241569
Rin118_2 in118_1 in118_2 9.241569
Rin118_3 in118_2 in118_3 9.241569
Rin118_4 in118_3 in118_4 9.241569
Rin118_5 in118_4 in118_5 9.241569
Rin118_6 in118_5 in118_6 9.241569
Rin118_7 in118_6 in118_7 9.241569
Rin118_8 in118_7 in118_8 9.241569
Rin118_9 in118_8 in118_9 9.241569
Rin118_10 in118_9 in118_10 9.241569
Rin118_11 in118_10 in118_11 9.241569
Rin118_12 in118_11 in118_12 9.241569
Rin118_13 in118_12 in118_13 9.241569
Rin118_14 in118_13 in118_14 9.241569
Rin118_15 in118_14 in118_15 9.241569
Rin118_16 in118_15 in118_16 9.241569
Rin118_17 in118_16 in118_17 9.241569
Rin118_18 in118_17 in118_18 9.241569
Rin118_19 in118_18 in118_19 9.241569
Rin118_20 in118_19 in118_20 9.241569
Rin118_21 in118_20 in118_21 9.241569
Rin118_22 in118_21 in118_22 9.241569
Rin118_23 in118_22 in118_23 9.241569
Rin118_24 in118_23 in118_24 9.241569
Rin118_25 in118_24 in118_25 9.241569
Rin118_26 in118_25 in118_26 9.241569
Rin118_27 in118_26 in118_27 9.241569
Rin118_28 in118_27 in118_28 9.241569
Rin118_29 in118 in118_29 9.241569
Rin118_30 in118_29 in118_30 9.241569
Rin118_31 in118_30 in118_31 9.241569
Rin118_32 in118_31 in118_32 9.241569
Rin118_33 in118_32 in118_33 9.241569
Rin118_34 in118_33 in118_34 9.241569
Rin118_35 in118_34 in118_35 9.241569
Rin118_36 in118_35 in118_36 9.241569
Rin118_37 in118_36 in118_37 9.241569
Rin118_38 in118_37 in118_38 9.241569
Rin118_39 in118_38 in118_39 9.241569
Rin118_40 in118_39 in118_40 9.241569
Rin118_41 in118_40 in118_41 9.241569
Rin118_42 in118_41 in118_42 9.241569
Rin118_43 in118_42 in118_43 9.241569
Rin118_44 in118_43 in118_44 9.241569
Rin118_45 in118_44 in118_45 9.241569
Rin118_46 in118_45 in118_46 9.241569
Rin118_47 in118_46 in118_47 9.241569
Rin118_48 in118_47 in118_48 9.241569
Rin118_49 in118_48 in118_49 9.241569
Rin118_50 in118_49 in118_50 9.241569
Rin118_51 in118_50 in118_51 9.241569
Rin118_52 in118_51 in118_52 9.241569
Rin118_53 in118_52 in118_53 9.241569
Rin118_54 in118_53 in118_54 9.241569
Rin118_55 in118_54 in118_55 9.241569
Rin118_56 in118_55 in118_56 9.241569
Rin118_57 in118 in118_57 9.241569
Rin118_58 in118_57 in118_58 9.241569
Rin118_59 in118_58 in118_59 9.241569
Rin118_60 in118_59 in118_60 9.241569
Rin118_61 in118_60 in118_61 9.241569
Rin118_62 in118_61 in118_62 9.241569
Rin118_63 in118_62 in118_63 9.241569
Rin118_64 in118_63 in118_64 9.241569
Rin118_65 in118_64 in118_65 9.241569
Rin118_66 in118_65 in118_66 9.241569
Rin118_67 in118_66 in118_67 9.241569
Rin118_68 in118_67 in118_68 9.241569
Rin118_69 in118_68 in118_69 9.241569
Rin118_70 in118_69 in118_70 9.241569
Rin118_71 in118_70 in118_71 9.241569
Rin118_72 in118_71 in118_72 9.241569
Rin118_73 in118_72 in118_73 9.241569
Rin118_74 in118_73 in118_74 9.241569
Rin118_75 in118_74 in118_75 9.241569
Rin118_76 in118_75 in118_76 9.241569
Rin118_77 in118_76 in118_77 9.241569
Rin118_78 in118_77 in118_78 9.241569
Rin118_79 in118_78 in118_79 9.241569
Rin118_80 in118_79 in118_80 9.241569
Rin118_81 in118_80 in118_81 9.241569
Rin118_82 in118_81 in118_82 9.241569
Rin118_83 in118_82 in118_83 9.241569
Rin118_84 in118_83 in118_84 9.241569
Rin119_1 in119 in119_1 9.241569
Rin119_2 in119_1 in119_2 9.241569
Rin119_3 in119_2 in119_3 9.241569
Rin119_4 in119_3 in119_4 9.241569
Rin119_5 in119_4 in119_5 9.241569
Rin119_6 in119_5 in119_6 9.241569
Rin119_7 in119_6 in119_7 9.241569
Rin119_8 in119_7 in119_8 9.241569
Rin119_9 in119_8 in119_9 9.241569
Rin119_10 in119_9 in119_10 9.241569
Rin119_11 in119_10 in119_11 9.241569
Rin119_12 in119_11 in119_12 9.241569
Rin119_13 in119_12 in119_13 9.241569
Rin119_14 in119_13 in119_14 9.241569
Rin119_15 in119_14 in119_15 9.241569
Rin119_16 in119_15 in119_16 9.241569
Rin119_17 in119_16 in119_17 9.241569
Rin119_18 in119_17 in119_18 9.241569
Rin119_19 in119_18 in119_19 9.241569
Rin119_20 in119_19 in119_20 9.241569
Rin119_21 in119_20 in119_21 9.241569
Rin119_22 in119_21 in119_22 9.241569
Rin119_23 in119_22 in119_23 9.241569
Rin119_24 in119_23 in119_24 9.241569
Rin119_25 in119_24 in119_25 9.241569
Rin119_26 in119_25 in119_26 9.241569
Rin119_27 in119_26 in119_27 9.241569
Rin119_28 in119_27 in119_28 9.241569
Rin119_29 in119 in119_29 9.241569
Rin119_30 in119_29 in119_30 9.241569
Rin119_31 in119_30 in119_31 9.241569
Rin119_32 in119_31 in119_32 9.241569
Rin119_33 in119_32 in119_33 9.241569
Rin119_34 in119_33 in119_34 9.241569
Rin119_35 in119_34 in119_35 9.241569
Rin119_36 in119_35 in119_36 9.241569
Rin119_37 in119_36 in119_37 9.241569
Rin119_38 in119_37 in119_38 9.241569
Rin119_39 in119_38 in119_39 9.241569
Rin119_40 in119_39 in119_40 9.241569
Rin119_41 in119_40 in119_41 9.241569
Rin119_42 in119_41 in119_42 9.241569
Rin119_43 in119_42 in119_43 9.241569
Rin119_44 in119_43 in119_44 9.241569
Rin119_45 in119_44 in119_45 9.241569
Rin119_46 in119_45 in119_46 9.241569
Rin119_47 in119_46 in119_47 9.241569
Rin119_48 in119_47 in119_48 9.241569
Rin119_49 in119_48 in119_49 9.241569
Rin119_50 in119_49 in119_50 9.241569
Rin119_51 in119_50 in119_51 9.241569
Rin119_52 in119_51 in119_52 9.241569
Rin119_53 in119_52 in119_53 9.241569
Rin119_54 in119_53 in119_54 9.241569
Rin119_55 in119_54 in119_55 9.241569
Rin119_56 in119_55 in119_56 9.241569
Rin119_57 in119 in119_57 9.241569
Rin119_58 in119_57 in119_58 9.241569
Rin119_59 in119_58 in119_59 9.241569
Rin119_60 in119_59 in119_60 9.241569
Rin119_61 in119_60 in119_61 9.241569
Rin119_62 in119_61 in119_62 9.241569
Rin119_63 in119_62 in119_63 9.241569
Rin119_64 in119_63 in119_64 9.241569
Rin119_65 in119_64 in119_65 9.241569
Rin119_66 in119_65 in119_66 9.241569
Rin119_67 in119_66 in119_67 9.241569
Rin119_68 in119_67 in119_68 9.241569
Rin119_69 in119_68 in119_69 9.241569
Rin119_70 in119_69 in119_70 9.241569
Rin119_71 in119_70 in119_71 9.241569
Rin119_72 in119_71 in119_72 9.241569
Rin119_73 in119_72 in119_73 9.241569
Rin119_74 in119_73 in119_74 9.241569
Rin119_75 in119_74 in119_75 9.241569
Rin119_76 in119_75 in119_76 9.241569
Rin119_77 in119_76 in119_77 9.241569
Rin119_78 in119_77 in119_78 9.241569
Rin119_79 in119_78 in119_79 9.241569
Rin119_80 in119_79 in119_80 9.241569
Rin119_81 in119_80 in119_81 9.241569
Rin119_82 in119_81 in119_82 9.241569
Rin119_83 in119_82 in119_83 9.241569
Rin119_84 in119_83 in119_84 9.241569
Rin120_1 in120 in120_1 9.241569
Rin120_2 in120_1 in120_2 9.241569
Rin120_3 in120_2 in120_3 9.241569
Rin120_4 in120_3 in120_4 9.241569
Rin120_5 in120_4 in120_5 9.241569
Rin120_6 in120_5 in120_6 9.241569
Rin120_7 in120_6 in120_7 9.241569
Rin120_8 in120_7 in120_8 9.241569
Rin120_9 in120_8 in120_9 9.241569
Rin120_10 in120_9 in120_10 9.241569
Rin120_11 in120_10 in120_11 9.241569
Rin120_12 in120_11 in120_12 9.241569
Rin120_13 in120_12 in120_13 9.241569
Rin120_14 in120_13 in120_14 9.241569
Rin120_15 in120_14 in120_15 9.241569
Rin120_16 in120_15 in120_16 9.241569
Rin120_17 in120_16 in120_17 9.241569
Rin120_18 in120_17 in120_18 9.241569
Rin120_19 in120_18 in120_19 9.241569
Rin120_20 in120_19 in120_20 9.241569
Rin120_21 in120_20 in120_21 9.241569
Rin120_22 in120_21 in120_22 9.241569
Rin120_23 in120_22 in120_23 9.241569
Rin120_24 in120_23 in120_24 9.241569
Rin120_25 in120_24 in120_25 9.241569
Rin120_26 in120_25 in120_26 9.241569
Rin120_27 in120_26 in120_27 9.241569
Rin120_28 in120_27 in120_28 9.241569
Rin120_29 in120 in120_29 9.241569
Rin120_30 in120_29 in120_30 9.241569
Rin120_31 in120_30 in120_31 9.241569
Rin120_32 in120_31 in120_32 9.241569
Rin120_33 in120_32 in120_33 9.241569
Rin120_34 in120_33 in120_34 9.241569
Rin120_35 in120_34 in120_35 9.241569
Rin120_36 in120_35 in120_36 9.241569
Rin120_37 in120_36 in120_37 9.241569
Rin120_38 in120_37 in120_38 9.241569
Rin120_39 in120_38 in120_39 9.241569
Rin120_40 in120_39 in120_40 9.241569
Rin120_41 in120_40 in120_41 9.241569
Rin120_42 in120_41 in120_42 9.241569
Rin120_43 in120_42 in120_43 9.241569
Rin120_44 in120_43 in120_44 9.241569
Rin120_45 in120_44 in120_45 9.241569
Rin120_46 in120_45 in120_46 9.241569
Rin120_47 in120_46 in120_47 9.241569
Rin120_48 in120_47 in120_48 9.241569
Rin120_49 in120_48 in120_49 9.241569
Rin120_50 in120_49 in120_50 9.241569
Rin120_51 in120_50 in120_51 9.241569
Rin120_52 in120_51 in120_52 9.241569
Rin120_53 in120_52 in120_53 9.241569
Rin120_54 in120_53 in120_54 9.241569
Rin120_55 in120_54 in120_55 9.241569
Rin120_56 in120_55 in120_56 9.241569
Rin120_57 in120 in120_57 9.241569
Rin120_58 in120_57 in120_58 9.241569
Rin120_59 in120_58 in120_59 9.241569
Rin120_60 in120_59 in120_60 9.241569
Rin120_61 in120_60 in120_61 9.241569
Rin120_62 in120_61 in120_62 9.241569
Rin120_63 in120_62 in120_63 9.241569
Rin120_64 in120_63 in120_64 9.241569
Rin120_65 in120_64 in120_65 9.241569
Rin120_66 in120_65 in120_66 9.241569
Rin120_67 in120_66 in120_67 9.241569
Rin120_68 in120_67 in120_68 9.241569
Rin120_69 in120_68 in120_69 9.241569
Rin120_70 in120_69 in120_70 9.241569
Rin120_71 in120_70 in120_71 9.241569
Rin120_72 in120_71 in120_72 9.241569
Rin120_73 in120_72 in120_73 9.241569
Rin120_74 in120_73 in120_74 9.241569
Rin120_75 in120_74 in120_75 9.241569
Rin120_76 in120_75 in120_76 9.241569
Rin120_77 in120_76 in120_77 9.241569
Rin120_78 in120_77 in120_78 9.241569
Rin120_79 in120_78 in120_79 9.241569
Rin120_80 in120_79 in120_80 9.241569
Rin120_81 in120_80 in120_81 9.241569
Rin120_82 in120_81 in120_82 9.241569
Rin120_83 in120_82 in120_83 9.241569
Rin120_84 in120_83 in120_84 9.241569
Rbias1 vdd vd1 9.241569
Rbias2 vd1 vd2 9.241569
Rbias3 vd2 vd3 9.241569
Rbias4 vd3 vd4 9.241569
Rbias5 vd4 vd5 9.241569
Rbias6 vd5 vd6 9.241569
Rbias7 vd6 vd7 9.241569
Rbias8 vd7 vd8 9.241569
Rbias9 vd8 vd9 9.241569
Rbias10 vd9 vd10 9.241569
Rbias11 vd10 vd11 9.241569
Rbias12 vd11 vd12 9.241569
Rbias13 vd12 vd13 9.241569
Rbias14 vd13 vd14 9.241569
Rbias15 vd14 vd15 9.241569
Rbias16 vd15 vd16 9.241569
Rbias17 vd16 vd17 9.241569
Rbias18 vd17 vd18 9.241569
Rbias19 vd18 vd19 9.241569
Rbias20 vd19 vd20 9.241569
Rbias21 vd20 vd21 9.241569
Rbias22 vd21 vd22 9.241569
Rbias23 vd22 vd23 9.241569
Rbias24 vd23 vd24 9.241569
Rbias25 vd24 vd25 9.241569
Rbias26 vd25 vd26 9.241569
Rbias27 vd26 vd27 9.241569
Rbias28 vd27 vd28 9.241569
Rbias29 vdd vd29 9.241569
Rbias30 vd29 vd30 9.241569
Rbias31 vd30 vd31 9.241569
Rbias32 vd31 vd32 9.241569
Rbias33 vd32 vd33 9.241569
Rbias34 vd33 vd34 9.241569
Rbias35 vd34 vd35 9.241569
Rbias36 vd35 vd36 9.241569
Rbias37 vd36 vd37 9.241569
Rbias38 vd37 vd38 9.241569
Rbias39 vd38 vd39 9.241569
Rbias40 vd39 vd40 9.241569
Rbias41 vd40 vd41 9.241569
Rbias42 vd41 vd42 9.241569
Rbias43 vd42 vd43 9.241569
Rbias44 vd43 vd44 9.241569
Rbias45 vd44 vd45 9.241569
Rbias46 vd45 vd46 9.241569
Rbias47 vd46 vd47 9.241569
Rbias48 vd47 vd48 9.241569
Rbias49 vd48 vd49 9.241569
Rbias50 vd49 vd50 9.241569
Rbias51 vd50 vd51 9.241569
Rbias52 vd51 vd52 9.241569
Rbias53 vd52 vd53 9.241569
Rbias54 vd53 vd54 9.241569
Rbias55 vd54 vd55 9.241569
Rbias56 vd55 vd56 9.241569
Rbias57 vdd vd57 9.241569
Rbias58 vd57 vd58 9.241569
Rbias59 vd58 vd59 9.241569
Rbias60 vd59 vd60 9.241569
Rbias61 vd60 vd61 9.241569
Rbias62 vd61 vd62 9.241569
Rbias63 vd62 vd63 9.241569
Rbias64 vd63 vd64 9.241569
Rbias65 vd64 vd65 9.241569
Rbias66 vd65 vd66 9.241569
Rbias67 vd66 vd67 9.241569
Rbias68 vd67 vd68 9.241569
Rbias69 vd68 vd69 9.241569
Rbias70 vd69 vd70 9.241569
Rbias71 vd70 vd71 9.241569
Rbias72 vd71 vd72 9.241569
Rbias73 vd72 vd73 9.241569
Rbias74 vd73 vd74 9.241569
Rbias75 vd74 vd75 9.241569
Rbias76 vd75 vd76 9.241569
Rbias77 vd76 vd77 9.241569
Rbias78 vd77 vd78 9.241569
Rbias79 vd78 vd79 9.241569
Rbias80 vd79 vd80 9.241569
Rbias81 vd80 vd81 9.241569
Rbias82 vd81 vd82 9.241569
Rbias83 vd82 vd83 9.241569
Rbias84 vd83 vd84 9.241569


**********Parasitic Resistances for I+ and I- Lines****************

Rsp1_1 sp1_1 sp2_1 11.551961
Rsn1_1 sn1_1 sn2_1 11.551961
Rsp1_2 sp1_2 sp2_2 11.551961
Rsn1_2 sn1_2 sn2_2 11.551961
Rsp1_3 sp1_3 sp2_3 11.551961
Rsn1_3 sn1_3 sn2_3 11.551961
Rsp1_4 sp1_4 sp2_4 11.551961
Rsn1_4 sn1_4 sn2_4 11.551961
Rsp1_5 sp1_5 sp2_5 11.551961
Rsn1_5 sn1_5 sn2_5 11.551961
Rsp1_6 sp1_6 sp2_6 11.551961
Rsn1_6 sn1_6 sn2_6 11.551961
Rsp1_7 sp1_7 sp2_7 11.551961
Rsn1_7 sn1_7 sn2_7 11.551961
Rsp1_8 sp1_8 sp2_8 11.551961
Rsn1_8 sn1_8 sn2_8 11.551961
Rsp1_9 sp1_9 sp2_9 11.551961
Rsn1_9 sn1_9 sn2_9 11.551961
Rsp1_10 sp1_10 sp2_10 11.551961
Rsn1_10 sn1_10 sn2_10 11.551961
Rsp1_11 sp1_11 sp2_11 11.551961
Rsn1_11 sn1_11 sn2_11 11.551961
Rsp1_12 sp1_12 sp2_12 11.551961
Rsn1_12 sn1_12 sn2_12 11.551961
Rsp1_13 sp1_13 sp2_13 11.551961
Rsn1_13 sn1_13 sn2_13 11.551961
Rsp1_14 sp1_14 sp2_14 11.551961
Rsn1_14 sn1_14 sn2_14 11.551961
Rsp1_15 sp1_15 sp2_15 11.551961
Rsn1_15 sn1_15 sn2_15 11.551961
Rsp1_16 sp1_16 sp2_16 11.551961
Rsn1_16 sn1_16 sn2_16 11.551961
Rsp1_17 sp1_17 sp2_17 11.551961
Rsn1_17 sn1_17 sn2_17 11.551961
Rsp1_18 sp1_18 sp2_18 11.551961
Rsn1_18 sn1_18 sn2_18 11.551961
Rsp1_19 sp1_19 sp2_19 11.551961
Rsn1_19 sn1_19 sn2_19 11.551961
Rsp1_20 sp1_20 sp2_20 11.551961
Rsn1_20 sn1_20 sn2_20 11.551961
Rsp1_21 sp1_21 sp2_21 11.551961
Rsn1_21 sn1_21 sn2_21 11.551961
Rsp1_22 sp1_22 sp2_22 11.551961
Rsn1_22 sn1_22 sn2_22 11.551961
Rsp1_23 sp1_23 sp2_23 11.551961
Rsn1_23 sn1_23 sn2_23 11.551961
Rsp1_24 sp1_24 sp2_24 11.551961
Rsn1_24 sn1_24 sn2_24 11.551961
Rsp1_25 sp1_25 sp2_25 11.551961
Rsn1_25 sn1_25 sn2_25 11.551961
Rsp1_26 sp1_26 sp2_26 11.551961
Rsn1_26 sn1_26 sn2_26 11.551961
Rsp1_27 sp1_27 sp2_27 11.551961
Rsn1_27 sn1_27 sn2_27 11.551961
Rsp1_28 sp1_28 sp2_28 11.551961
Rsn1_28 sn1_28 sn2_28 11.551961
Rsp1_29 sp1_29 sp2_29 11.551961
Rsn1_29 sn1_29 sn2_29 11.551961
Rsp1_30 sp1_30 sp2_30 11.551961
Rsn1_30 sn1_30 sn2_30 11.551961
Rsp1_31 sp1_31 sp2_31 11.551961
Rsn1_31 sn1_31 sn2_31 11.551961
Rsp1_32 sp1_32 sp2_32 11.551961
Rsn1_32 sn1_32 sn2_32 11.551961
Rsp1_33 sp1_33 sp2_33 11.551961
Rsn1_33 sn1_33 sn2_33 11.551961
Rsp1_34 sp1_34 sp2_34 11.551961
Rsn1_34 sn1_34 sn2_34 11.551961
Rsp1_35 sp1_35 sp2_35 11.551961
Rsn1_35 sn1_35 sn2_35 11.551961
Rsp1_36 sp1_36 sp2_36 11.551961
Rsn1_36 sn1_36 sn2_36 11.551961
Rsp1_37 sp1_37 sp2_37 11.551961
Rsn1_37 sn1_37 sn2_37 11.551961
Rsp1_38 sp1_38 sp2_38 11.551961
Rsn1_38 sn1_38 sn2_38 11.551961
Rsp1_39 sp1_39 sp2_39 11.551961
Rsn1_39 sn1_39 sn2_39 11.551961
Rsp1_40 sp1_40 sp2_40 11.551961
Rsn1_40 sn1_40 sn2_40 11.551961
Rsp1_41 sp1_41 sp2_41 11.551961
Rsn1_41 sn1_41 sn2_41 11.551961
Rsp1_42 sp1_42 sp2_42 11.551961
Rsn1_42 sn1_42 sn2_42 11.551961
Rsp1_43 sp1_43 sp2_43 11.551961
Rsn1_43 sn1_43 sn2_43 11.551961
Rsp1_44 sp1_44 sp2_44 11.551961
Rsn1_44 sn1_44 sn2_44 11.551961
Rsp1_45 sp1_45 sp2_45 11.551961
Rsn1_45 sn1_45 sn2_45 11.551961
Rsp1_46 sp1_46 sp2_46 11.551961
Rsn1_46 sn1_46 sn2_46 11.551961
Rsp1_47 sp1_47 sp2_47 11.551961
Rsn1_47 sn1_47 sn2_47 11.551961
Rsp1_48 sp1_48 sp2_48 11.551961
Rsn1_48 sn1_48 sn2_48 11.551961
Rsp1_49 sp1_49 sp2_49 11.551961
Rsn1_49 sn1_49 sn2_49 11.551961
Rsp1_50 sp1_50 sp2_50 11.551961
Rsn1_50 sn1_50 sn2_50 11.551961
Rsp1_51 sp1_51 sp2_51 11.551961
Rsn1_51 sn1_51 sn2_51 11.551961
Rsp1_52 sp1_52 sp2_52 11.551961
Rsn1_52 sn1_52 sn2_52 11.551961
Rsp1_53 sp1_53 sp2_53 11.551961
Rsn1_53 sn1_53 sn2_53 11.551961
Rsp1_54 sp1_54 sp2_54 11.551961
Rsn1_54 sn1_54 sn2_54 11.551961
Rsp1_55 sp1_55 sp2_55 11.551961
Rsn1_55 sn1_55 sn2_55 11.551961
Rsp1_56 sp1_56 sp2_56 11.551961
Rsn1_56 sn1_56 sn2_56 11.551961
Rsp1_57 sp1_57 sp2_57 11.551961
Rsn1_57 sn1_57 sn2_57 11.551961
Rsp1_58 sp1_58 sp2_58 11.551961
Rsn1_58 sn1_58 sn2_58 11.551961
Rsp1_59 sp1_59 sp2_59 11.551961
Rsn1_59 sn1_59 sn2_59 11.551961
Rsp1_60 sp1_60 sp2_60 11.551961
Rsn1_60 sn1_60 sn2_60 11.551961
Rsp1_61 sp1_61 sp2_61 11.551961
Rsn1_61 sn1_61 sn2_61 11.551961
Rsp1_62 sp1_62 sp2_62 11.551961
Rsn1_62 sn1_62 sn2_62 11.551961
Rsp1_63 sp1_63 sp2_63 11.551961
Rsn1_63 sn1_63 sn2_63 11.551961
Rsp1_64 sp1_64 sp2_64 11.551961
Rsn1_64 sn1_64 sn2_64 11.551961
Rsp1_65 sp1_65 sp2_65 11.551961
Rsn1_65 sn1_65 sn2_65 11.551961
Rsp1_66 sp1_66 sp2_66 11.551961
Rsn1_66 sn1_66 sn2_66 11.551961
Rsp1_67 sp1_67 sp2_67 11.551961
Rsn1_67 sn1_67 sn2_67 11.551961
Rsp1_68 sp1_68 sp2_68 11.551961
Rsn1_68 sn1_68 sn2_68 11.551961
Rsp1_69 sp1_69 sp2_69 11.551961
Rsn1_69 sn1_69 sn2_69 11.551961
Rsp1_70 sp1_70 sp2_70 11.551961
Rsn1_70 sn1_70 sn2_70 11.551961
Rsp1_71 sp1_71 sp2_71 11.551961
Rsn1_71 sn1_71 sn2_71 11.551961
Rsp1_72 sp1_72 sp2_72 11.551961
Rsn1_72 sn1_72 sn2_72 11.551961
Rsp1_73 sp1_73 sp2_73 11.551961
Rsn1_73 sn1_73 sn2_73 11.551961
Rsp1_74 sp1_74 sp2_74 11.551961
Rsn1_74 sn1_74 sn2_74 11.551961
Rsp1_75 sp1_75 sp2_75 11.551961
Rsn1_75 sn1_75 sn2_75 11.551961
Rsp1_76 sp1_76 sp2_76 11.551961
Rsn1_76 sn1_76 sn2_76 11.551961
Rsp1_77 sp1_77 sp2_77 11.551961
Rsn1_77 sn1_77 sn2_77 11.551961
Rsp1_78 sp1_78 sp2_78 11.551961
Rsn1_78 sn1_78 sn2_78 11.551961
Rsp1_79 sp1_79 sp2_79 11.551961
Rsn1_79 sn1_79 sn2_79 11.551961
Rsp1_80 sp1_80 sp2_80 11.551961
Rsn1_80 sn1_80 sn2_80 11.551961
Rsp1_81 sp1_81 sp2_81 11.551961
Rsn1_81 sn1_81 sn2_81 11.551961
Rsp1_82 sp1_82 sp2_82 11.551961
Rsn1_82 sn1_82 sn2_82 11.551961
Rsp1_83 sp1_83 sp2_83 11.551961
Rsn1_83 sn1_83 sn2_83 11.551961
Rsp1_84 sp1_84 sp2_84 11.551961
Rsn1_84 sn1_84 sn2_84 11.551961
Rsp2_1 sp2_1 sp3_1 11.551961
Rsn2_1 sn2_1 sn3_1 11.551961
Rsp2_2 sp2_2 sp3_2 11.551961
Rsn2_2 sn2_2 sn3_2 11.551961
Rsp2_3 sp2_3 sp3_3 11.551961
Rsn2_3 sn2_3 sn3_3 11.551961
Rsp2_4 sp2_4 sp3_4 11.551961
Rsn2_4 sn2_4 sn3_4 11.551961
Rsp2_5 sp2_5 sp3_5 11.551961
Rsn2_5 sn2_5 sn3_5 11.551961
Rsp2_6 sp2_6 sp3_6 11.551961
Rsn2_6 sn2_6 sn3_6 11.551961
Rsp2_7 sp2_7 sp3_7 11.551961
Rsn2_7 sn2_7 sn3_7 11.551961
Rsp2_8 sp2_8 sp3_8 11.551961
Rsn2_8 sn2_8 sn3_8 11.551961
Rsp2_9 sp2_9 sp3_9 11.551961
Rsn2_9 sn2_9 sn3_9 11.551961
Rsp2_10 sp2_10 sp3_10 11.551961
Rsn2_10 sn2_10 sn3_10 11.551961
Rsp2_11 sp2_11 sp3_11 11.551961
Rsn2_11 sn2_11 sn3_11 11.551961
Rsp2_12 sp2_12 sp3_12 11.551961
Rsn2_12 sn2_12 sn3_12 11.551961
Rsp2_13 sp2_13 sp3_13 11.551961
Rsn2_13 sn2_13 sn3_13 11.551961
Rsp2_14 sp2_14 sp3_14 11.551961
Rsn2_14 sn2_14 sn3_14 11.551961
Rsp2_15 sp2_15 sp3_15 11.551961
Rsn2_15 sn2_15 sn3_15 11.551961
Rsp2_16 sp2_16 sp3_16 11.551961
Rsn2_16 sn2_16 sn3_16 11.551961
Rsp2_17 sp2_17 sp3_17 11.551961
Rsn2_17 sn2_17 sn3_17 11.551961
Rsp2_18 sp2_18 sp3_18 11.551961
Rsn2_18 sn2_18 sn3_18 11.551961
Rsp2_19 sp2_19 sp3_19 11.551961
Rsn2_19 sn2_19 sn3_19 11.551961
Rsp2_20 sp2_20 sp3_20 11.551961
Rsn2_20 sn2_20 sn3_20 11.551961
Rsp2_21 sp2_21 sp3_21 11.551961
Rsn2_21 sn2_21 sn3_21 11.551961
Rsp2_22 sp2_22 sp3_22 11.551961
Rsn2_22 sn2_22 sn3_22 11.551961
Rsp2_23 sp2_23 sp3_23 11.551961
Rsn2_23 sn2_23 sn3_23 11.551961
Rsp2_24 sp2_24 sp3_24 11.551961
Rsn2_24 sn2_24 sn3_24 11.551961
Rsp2_25 sp2_25 sp3_25 11.551961
Rsn2_25 sn2_25 sn3_25 11.551961
Rsp2_26 sp2_26 sp3_26 11.551961
Rsn2_26 sn2_26 sn3_26 11.551961
Rsp2_27 sp2_27 sp3_27 11.551961
Rsn2_27 sn2_27 sn3_27 11.551961
Rsp2_28 sp2_28 sp3_28 11.551961
Rsn2_28 sn2_28 sn3_28 11.551961
Rsp2_29 sp2_29 sp3_29 11.551961
Rsn2_29 sn2_29 sn3_29 11.551961
Rsp2_30 sp2_30 sp3_30 11.551961
Rsn2_30 sn2_30 sn3_30 11.551961
Rsp2_31 sp2_31 sp3_31 11.551961
Rsn2_31 sn2_31 sn3_31 11.551961
Rsp2_32 sp2_32 sp3_32 11.551961
Rsn2_32 sn2_32 sn3_32 11.551961
Rsp2_33 sp2_33 sp3_33 11.551961
Rsn2_33 sn2_33 sn3_33 11.551961
Rsp2_34 sp2_34 sp3_34 11.551961
Rsn2_34 sn2_34 sn3_34 11.551961
Rsp2_35 sp2_35 sp3_35 11.551961
Rsn2_35 sn2_35 sn3_35 11.551961
Rsp2_36 sp2_36 sp3_36 11.551961
Rsn2_36 sn2_36 sn3_36 11.551961
Rsp2_37 sp2_37 sp3_37 11.551961
Rsn2_37 sn2_37 sn3_37 11.551961
Rsp2_38 sp2_38 sp3_38 11.551961
Rsn2_38 sn2_38 sn3_38 11.551961
Rsp2_39 sp2_39 sp3_39 11.551961
Rsn2_39 sn2_39 sn3_39 11.551961
Rsp2_40 sp2_40 sp3_40 11.551961
Rsn2_40 sn2_40 sn3_40 11.551961
Rsp2_41 sp2_41 sp3_41 11.551961
Rsn2_41 sn2_41 sn3_41 11.551961
Rsp2_42 sp2_42 sp3_42 11.551961
Rsn2_42 sn2_42 sn3_42 11.551961
Rsp2_43 sp2_43 sp3_43 11.551961
Rsn2_43 sn2_43 sn3_43 11.551961
Rsp2_44 sp2_44 sp3_44 11.551961
Rsn2_44 sn2_44 sn3_44 11.551961
Rsp2_45 sp2_45 sp3_45 11.551961
Rsn2_45 sn2_45 sn3_45 11.551961
Rsp2_46 sp2_46 sp3_46 11.551961
Rsn2_46 sn2_46 sn3_46 11.551961
Rsp2_47 sp2_47 sp3_47 11.551961
Rsn2_47 sn2_47 sn3_47 11.551961
Rsp2_48 sp2_48 sp3_48 11.551961
Rsn2_48 sn2_48 sn3_48 11.551961
Rsp2_49 sp2_49 sp3_49 11.551961
Rsn2_49 sn2_49 sn3_49 11.551961
Rsp2_50 sp2_50 sp3_50 11.551961
Rsn2_50 sn2_50 sn3_50 11.551961
Rsp2_51 sp2_51 sp3_51 11.551961
Rsn2_51 sn2_51 sn3_51 11.551961
Rsp2_52 sp2_52 sp3_52 11.551961
Rsn2_52 sn2_52 sn3_52 11.551961
Rsp2_53 sp2_53 sp3_53 11.551961
Rsn2_53 sn2_53 sn3_53 11.551961
Rsp2_54 sp2_54 sp3_54 11.551961
Rsn2_54 sn2_54 sn3_54 11.551961
Rsp2_55 sp2_55 sp3_55 11.551961
Rsn2_55 sn2_55 sn3_55 11.551961
Rsp2_56 sp2_56 sp3_56 11.551961
Rsn2_56 sn2_56 sn3_56 11.551961
Rsp2_57 sp2_57 sp3_57 11.551961
Rsn2_57 sn2_57 sn3_57 11.551961
Rsp2_58 sp2_58 sp3_58 11.551961
Rsn2_58 sn2_58 sn3_58 11.551961
Rsp2_59 sp2_59 sp3_59 11.551961
Rsn2_59 sn2_59 sn3_59 11.551961
Rsp2_60 sp2_60 sp3_60 11.551961
Rsn2_60 sn2_60 sn3_60 11.551961
Rsp2_61 sp2_61 sp3_61 11.551961
Rsn2_61 sn2_61 sn3_61 11.551961
Rsp2_62 sp2_62 sp3_62 11.551961
Rsn2_62 sn2_62 sn3_62 11.551961
Rsp2_63 sp2_63 sp3_63 11.551961
Rsn2_63 sn2_63 sn3_63 11.551961
Rsp2_64 sp2_64 sp3_64 11.551961
Rsn2_64 sn2_64 sn3_64 11.551961
Rsp2_65 sp2_65 sp3_65 11.551961
Rsn2_65 sn2_65 sn3_65 11.551961
Rsp2_66 sp2_66 sp3_66 11.551961
Rsn2_66 sn2_66 sn3_66 11.551961
Rsp2_67 sp2_67 sp3_67 11.551961
Rsn2_67 sn2_67 sn3_67 11.551961
Rsp2_68 sp2_68 sp3_68 11.551961
Rsn2_68 sn2_68 sn3_68 11.551961
Rsp2_69 sp2_69 sp3_69 11.551961
Rsn2_69 sn2_69 sn3_69 11.551961
Rsp2_70 sp2_70 sp3_70 11.551961
Rsn2_70 sn2_70 sn3_70 11.551961
Rsp2_71 sp2_71 sp3_71 11.551961
Rsn2_71 sn2_71 sn3_71 11.551961
Rsp2_72 sp2_72 sp3_72 11.551961
Rsn2_72 sn2_72 sn3_72 11.551961
Rsp2_73 sp2_73 sp3_73 11.551961
Rsn2_73 sn2_73 sn3_73 11.551961
Rsp2_74 sp2_74 sp3_74 11.551961
Rsn2_74 sn2_74 sn3_74 11.551961
Rsp2_75 sp2_75 sp3_75 11.551961
Rsn2_75 sn2_75 sn3_75 11.551961
Rsp2_76 sp2_76 sp3_76 11.551961
Rsn2_76 sn2_76 sn3_76 11.551961
Rsp2_77 sp2_77 sp3_77 11.551961
Rsn2_77 sn2_77 sn3_77 11.551961
Rsp2_78 sp2_78 sp3_78 11.551961
Rsn2_78 sn2_78 sn3_78 11.551961
Rsp2_79 sp2_79 sp3_79 11.551961
Rsn2_79 sn2_79 sn3_79 11.551961
Rsp2_80 sp2_80 sp3_80 11.551961
Rsn2_80 sn2_80 sn3_80 11.551961
Rsp2_81 sp2_81 sp3_81 11.551961
Rsn2_81 sn2_81 sn3_81 11.551961
Rsp2_82 sp2_82 sp3_82 11.551961
Rsn2_82 sn2_82 sn3_82 11.551961
Rsp2_83 sp2_83 sp3_83 11.551961
Rsn2_83 sn2_83 sn3_83 11.551961
Rsp2_84 sp2_84 sp3_84 11.551961
Rsn2_84 sn2_84 sn3_84 11.551961
Rsp3_1 sp3_1 sp4_1 11.551961
Rsn3_1 sn3_1 sn4_1 11.551961
Rsp3_2 sp3_2 sp4_2 11.551961
Rsn3_2 sn3_2 sn4_2 11.551961
Rsp3_3 sp3_3 sp4_3 11.551961
Rsn3_3 sn3_3 sn4_3 11.551961
Rsp3_4 sp3_4 sp4_4 11.551961
Rsn3_4 sn3_4 sn4_4 11.551961
Rsp3_5 sp3_5 sp4_5 11.551961
Rsn3_5 sn3_5 sn4_5 11.551961
Rsp3_6 sp3_6 sp4_6 11.551961
Rsn3_6 sn3_6 sn4_6 11.551961
Rsp3_7 sp3_7 sp4_7 11.551961
Rsn3_7 sn3_7 sn4_7 11.551961
Rsp3_8 sp3_8 sp4_8 11.551961
Rsn3_8 sn3_8 sn4_8 11.551961
Rsp3_9 sp3_9 sp4_9 11.551961
Rsn3_9 sn3_9 sn4_9 11.551961
Rsp3_10 sp3_10 sp4_10 11.551961
Rsn3_10 sn3_10 sn4_10 11.551961
Rsp3_11 sp3_11 sp4_11 11.551961
Rsn3_11 sn3_11 sn4_11 11.551961
Rsp3_12 sp3_12 sp4_12 11.551961
Rsn3_12 sn3_12 sn4_12 11.551961
Rsp3_13 sp3_13 sp4_13 11.551961
Rsn3_13 sn3_13 sn4_13 11.551961
Rsp3_14 sp3_14 sp4_14 11.551961
Rsn3_14 sn3_14 sn4_14 11.551961
Rsp3_15 sp3_15 sp4_15 11.551961
Rsn3_15 sn3_15 sn4_15 11.551961
Rsp3_16 sp3_16 sp4_16 11.551961
Rsn3_16 sn3_16 sn4_16 11.551961
Rsp3_17 sp3_17 sp4_17 11.551961
Rsn3_17 sn3_17 sn4_17 11.551961
Rsp3_18 sp3_18 sp4_18 11.551961
Rsn3_18 sn3_18 sn4_18 11.551961
Rsp3_19 sp3_19 sp4_19 11.551961
Rsn3_19 sn3_19 sn4_19 11.551961
Rsp3_20 sp3_20 sp4_20 11.551961
Rsn3_20 sn3_20 sn4_20 11.551961
Rsp3_21 sp3_21 sp4_21 11.551961
Rsn3_21 sn3_21 sn4_21 11.551961
Rsp3_22 sp3_22 sp4_22 11.551961
Rsn3_22 sn3_22 sn4_22 11.551961
Rsp3_23 sp3_23 sp4_23 11.551961
Rsn3_23 sn3_23 sn4_23 11.551961
Rsp3_24 sp3_24 sp4_24 11.551961
Rsn3_24 sn3_24 sn4_24 11.551961
Rsp3_25 sp3_25 sp4_25 11.551961
Rsn3_25 sn3_25 sn4_25 11.551961
Rsp3_26 sp3_26 sp4_26 11.551961
Rsn3_26 sn3_26 sn4_26 11.551961
Rsp3_27 sp3_27 sp4_27 11.551961
Rsn3_27 sn3_27 sn4_27 11.551961
Rsp3_28 sp3_28 sp4_28 11.551961
Rsn3_28 sn3_28 sn4_28 11.551961
Rsp3_29 sp3_29 sp4_29 11.551961
Rsn3_29 sn3_29 sn4_29 11.551961
Rsp3_30 sp3_30 sp4_30 11.551961
Rsn3_30 sn3_30 sn4_30 11.551961
Rsp3_31 sp3_31 sp4_31 11.551961
Rsn3_31 sn3_31 sn4_31 11.551961
Rsp3_32 sp3_32 sp4_32 11.551961
Rsn3_32 sn3_32 sn4_32 11.551961
Rsp3_33 sp3_33 sp4_33 11.551961
Rsn3_33 sn3_33 sn4_33 11.551961
Rsp3_34 sp3_34 sp4_34 11.551961
Rsn3_34 sn3_34 sn4_34 11.551961
Rsp3_35 sp3_35 sp4_35 11.551961
Rsn3_35 sn3_35 sn4_35 11.551961
Rsp3_36 sp3_36 sp4_36 11.551961
Rsn3_36 sn3_36 sn4_36 11.551961
Rsp3_37 sp3_37 sp4_37 11.551961
Rsn3_37 sn3_37 sn4_37 11.551961
Rsp3_38 sp3_38 sp4_38 11.551961
Rsn3_38 sn3_38 sn4_38 11.551961
Rsp3_39 sp3_39 sp4_39 11.551961
Rsn3_39 sn3_39 sn4_39 11.551961
Rsp3_40 sp3_40 sp4_40 11.551961
Rsn3_40 sn3_40 sn4_40 11.551961
Rsp3_41 sp3_41 sp4_41 11.551961
Rsn3_41 sn3_41 sn4_41 11.551961
Rsp3_42 sp3_42 sp4_42 11.551961
Rsn3_42 sn3_42 sn4_42 11.551961
Rsp3_43 sp3_43 sp4_43 11.551961
Rsn3_43 sn3_43 sn4_43 11.551961
Rsp3_44 sp3_44 sp4_44 11.551961
Rsn3_44 sn3_44 sn4_44 11.551961
Rsp3_45 sp3_45 sp4_45 11.551961
Rsn3_45 sn3_45 sn4_45 11.551961
Rsp3_46 sp3_46 sp4_46 11.551961
Rsn3_46 sn3_46 sn4_46 11.551961
Rsp3_47 sp3_47 sp4_47 11.551961
Rsn3_47 sn3_47 sn4_47 11.551961
Rsp3_48 sp3_48 sp4_48 11.551961
Rsn3_48 sn3_48 sn4_48 11.551961
Rsp3_49 sp3_49 sp4_49 11.551961
Rsn3_49 sn3_49 sn4_49 11.551961
Rsp3_50 sp3_50 sp4_50 11.551961
Rsn3_50 sn3_50 sn4_50 11.551961
Rsp3_51 sp3_51 sp4_51 11.551961
Rsn3_51 sn3_51 sn4_51 11.551961
Rsp3_52 sp3_52 sp4_52 11.551961
Rsn3_52 sn3_52 sn4_52 11.551961
Rsp3_53 sp3_53 sp4_53 11.551961
Rsn3_53 sn3_53 sn4_53 11.551961
Rsp3_54 sp3_54 sp4_54 11.551961
Rsn3_54 sn3_54 sn4_54 11.551961
Rsp3_55 sp3_55 sp4_55 11.551961
Rsn3_55 sn3_55 sn4_55 11.551961
Rsp3_56 sp3_56 sp4_56 11.551961
Rsn3_56 sn3_56 sn4_56 11.551961
Rsp3_57 sp3_57 sp4_57 11.551961
Rsn3_57 sn3_57 sn4_57 11.551961
Rsp3_58 sp3_58 sp4_58 11.551961
Rsn3_58 sn3_58 sn4_58 11.551961
Rsp3_59 sp3_59 sp4_59 11.551961
Rsn3_59 sn3_59 sn4_59 11.551961
Rsp3_60 sp3_60 sp4_60 11.551961
Rsn3_60 sn3_60 sn4_60 11.551961
Rsp3_61 sp3_61 sp4_61 11.551961
Rsn3_61 sn3_61 sn4_61 11.551961
Rsp3_62 sp3_62 sp4_62 11.551961
Rsn3_62 sn3_62 sn4_62 11.551961
Rsp3_63 sp3_63 sp4_63 11.551961
Rsn3_63 sn3_63 sn4_63 11.551961
Rsp3_64 sp3_64 sp4_64 11.551961
Rsn3_64 sn3_64 sn4_64 11.551961
Rsp3_65 sp3_65 sp4_65 11.551961
Rsn3_65 sn3_65 sn4_65 11.551961
Rsp3_66 sp3_66 sp4_66 11.551961
Rsn3_66 sn3_66 sn4_66 11.551961
Rsp3_67 sp3_67 sp4_67 11.551961
Rsn3_67 sn3_67 sn4_67 11.551961
Rsp3_68 sp3_68 sp4_68 11.551961
Rsn3_68 sn3_68 sn4_68 11.551961
Rsp3_69 sp3_69 sp4_69 11.551961
Rsn3_69 sn3_69 sn4_69 11.551961
Rsp3_70 sp3_70 sp4_70 11.551961
Rsn3_70 sn3_70 sn4_70 11.551961
Rsp3_71 sp3_71 sp4_71 11.551961
Rsn3_71 sn3_71 sn4_71 11.551961
Rsp3_72 sp3_72 sp4_72 11.551961
Rsn3_72 sn3_72 sn4_72 11.551961
Rsp3_73 sp3_73 sp4_73 11.551961
Rsn3_73 sn3_73 sn4_73 11.551961
Rsp3_74 sp3_74 sp4_74 11.551961
Rsn3_74 sn3_74 sn4_74 11.551961
Rsp3_75 sp3_75 sp4_75 11.551961
Rsn3_75 sn3_75 sn4_75 11.551961
Rsp3_76 sp3_76 sp4_76 11.551961
Rsn3_76 sn3_76 sn4_76 11.551961
Rsp3_77 sp3_77 sp4_77 11.551961
Rsn3_77 sn3_77 sn4_77 11.551961
Rsp3_78 sp3_78 sp4_78 11.551961
Rsn3_78 sn3_78 sn4_78 11.551961
Rsp3_79 sp3_79 sp4_79 11.551961
Rsn3_79 sn3_79 sn4_79 11.551961
Rsp3_80 sp3_80 sp4_80 11.551961
Rsn3_80 sn3_80 sn4_80 11.551961
Rsp3_81 sp3_81 sp4_81 11.551961
Rsn3_81 sn3_81 sn4_81 11.551961
Rsp3_82 sp3_82 sp4_82 11.551961
Rsn3_82 sn3_82 sn4_82 11.551961
Rsp3_83 sp3_83 sp4_83 11.551961
Rsn3_83 sn3_83 sn4_83 11.551961
Rsp3_84 sp3_84 sp4_84 11.551961
Rsn3_84 sn3_84 sn4_84 11.551961
Rsp4_1 sp4_1 sp5_1 11.551961
Rsn4_1 sn4_1 sn5_1 11.551961
Rsp4_2 sp4_2 sp5_2 11.551961
Rsn4_2 sn4_2 sn5_2 11.551961
Rsp4_3 sp4_3 sp5_3 11.551961
Rsn4_3 sn4_3 sn5_3 11.551961
Rsp4_4 sp4_4 sp5_4 11.551961
Rsn4_4 sn4_4 sn5_4 11.551961
Rsp4_5 sp4_5 sp5_5 11.551961
Rsn4_5 sn4_5 sn5_5 11.551961
Rsp4_6 sp4_6 sp5_6 11.551961
Rsn4_6 sn4_6 sn5_6 11.551961
Rsp4_7 sp4_7 sp5_7 11.551961
Rsn4_7 sn4_7 sn5_7 11.551961
Rsp4_8 sp4_8 sp5_8 11.551961
Rsn4_8 sn4_8 sn5_8 11.551961
Rsp4_9 sp4_9 sp5_9 11.551961
Rsn4_9 sn4_9 sn5_9 11.551961
Rsp4_10 sp4_10 sp5_10 11.551961
Rsn4_10 sn4_10 sn5_10 11.551961
Rsp4_11 sp4_11 sp5_11 11.551961
Rsn4_11 sn4_11 sn5_11 11.551961
Rsp4_12 sp4_12 sp5_12 11.551961
Rsn4_12 sn4_12 sn5_12 11.551961
Rsp4_13 sp4_13 sp5_13 11.551961
Rsn4_13 sn4_13 sn5_13 11.551961
Rsp4_14 sp4_14 sp5_14 11.551961
Rsn4_14 sn4_14 sn5_14 11.551961
Rsp4_15 sp4_15 sp5_15 11.551961
Rsn4_15 sn4_15 sn5_15 11.551961
Rsp4_16 sp4_16 sp5_16 11.551961
Rsn4_16 sn4_16 sn5_16 11.551961
Rsp4_17 sp4_17 sp5_17 11.551961
Rsn4_17 sn4_17 sn5_17 11.551961
Rsp4_18 sp4_18 sp5_18 11.551961
Rsn4_18 sn4_18 sn5_18 11.551961
Rsp4_19 sp4_19 sp5_19 11.551961
Rsn4_19 sn4_19 sn5_19 11.551961
Rsp4_20 sp4_20 sp5_20 11.551961
Rsn4_20 sn4_20 sn5_20 11.551961
Rsp4_21 sp4_21 sp5_21 11.551961
Rsn4_21 sn4_21 sn5_21 11.551961
Rsp4_22 sp4_22 sp5_22 11.551961
Rsn4_22 sn4_22 sn5_22 11.551961
Rsp4_23 sp4_23 sp5_23 11.551961
Rsn4_23 sn4_23 sn5_23 11.551961
Rsp4_24 sp4_24 sp5_24 11.551961
Rsn4_24 sn4_24 sn5_24 11.551961
Rsp4_25 sp4_25 sp5_25 11.551961
Rsn4_25 sn4_25 sn5_25 11.551961
Rsp4_26 sp4_26 sp5_26 11.551961
Rsn4_26 sn4_26 sn5_26 11.551961
Rsp4_27 sp4_27 sp5_27 11.551961
Rsn4_27 sn4_27 sn5_27 11.551961
Rsp4_28 sp4_28 sp5_28 11.551961
Rsn4_28 sn4_28 sn5_28 11.551961
Rsp4_29 sp4_29 sp5_29 11.551961
Rsn4_29 sn4_29 sn5_29 11.551961
Rsp4_30 sp4_30 sp5_30 11.551961
Rsn4_30 sn4_30 sn5_30 11.551961
Rsp4_31 sp4_31 sp5_31 11.551961
Rsn4_31 sn4_31 sn5_31 11.551961
Rsp4_32 sp4_32 sp5_32 11.551961
Rsn4_32 sn4_32 sn5_32 11.551961
Rsp4_33 sp4_33 sp5_33 11.551961
Rsn4_33 sn4_33 sn5_33 11.551961
Rsp4_34 sp4_34 sp5_34 11.551961
Rsn4_34 sn4_34 sn5_34 11.551961
Rsp4_35 sp4_35 sp5_35 11.551961
Rsn4_35 sn4_35 sn5_35 11.551961
Rsp4_36 sp4_36 sp5_36 11.551961
Rsn4_36 sn4_36 sn5_36 11.551961
Rsp4_37 sp4_37 sp5_37 11.551961
Rsn4_37 sn4_37 sn5_37 11.551961
Rsp4_38 sp4_38 sp5_38 11.551961
Rsn4_38 sn4_38 sn5_38 11.551961
Rsp4_39 sp4_39 sp5_39 11.551961
Rsn4_39 sn4_39 sn5_39 11.551961
Rsp4_40 sp4_40 sp5_40 11.551961
Rsn4_40 sn4_40 sn5_40 11.551961
Rsp4_41 sp4_41 sp5_41 11.551961
Rsn4_41 sn4_41 sn5_41 11.551961
Rsp4_42 sp4_42 sp5_42 11.551961
Rsn4_42 sn4_42 sn5_42 11.551961
Rsp4_43 sp4_43 sp5_43 11.551961
Rsn4_43 sn4_43 sn5_43 11.551961
Rsp4_44 sp4_44 sp5_44 11.551961
Rsn4_44 sn4_44 sn5_44 11.551961
Rsp4_45 sp4_45 sp5_45 11.551961
Rsn4_45 sn4_45 sn5_45 11.551961
Rsp4_46 sp4_46 sp5_46 11.551961
Rsn4_46 sn4_46 sn5_46 11.551961
Rsp4_47 sp4_47 sp5_47 11.551961
Rsn4_47 sn4_47 sn5_47 11.551961
Rsp4_48 sp4_48 sp5_48 11.551961
Rsn4_48 sn4_48 sn5_48 11.551961
Rsp4_49 sp4_49 sp5_49 11.551961
Rsn4_49 sn4_49 sn5_49 11.551961
Rsp4_50 sp4_50 sp5_50 11.551961
Rsn4_50 sn4_50 sn5_50 11.551961
Rsp4_51 sp4_51 sp5_51 11.551961
Rsn4_51 sn4_51 sn5_51 11.551961
Rsp4_52 sp4_52 sp5_52 11.551961
Rsn4_52 sn4_52 sn5_52 11.551961
Rsp4_53 sp4_53 sp5_53 11.551961
Rsn4_53 sn4_53 sn5_53 11.551961
Rsp4_54 sp4_54 sp5_54 11.551961
Rsn4_54 sn4_54 sn5_54 11.551961
Rsp4_55 sp4_55 sp5_55 11.551961
Rsn4_55 sn4_55 sn5_55 11.551961
Rsp4_56 sp4_56 sp5_56 11.551961
Rsn4_56 sn4_56 sn5_56 11.551961
Rsp4_57 sp4_57 sp5_57 11.551961
Rsn4_57 sn4_57 sn5_57 11.551961
Rsp4_58 sp4_58 sp5_58 11.551961
Rsn4_58 sn4_58 sn5_58 11.551961
Rsp4_59 sp4_59 sp5_59 11.551961
Rsn4_59 sn4_59 sn5_59 11.551961
Rsp4_60 sp4_60 sp5_60 11.551961
Rsn4_60 sn4_60 sn5_60 11.551961
Rsp4_61 sp4_61 sp5_61 11.551961
Rsn4_61 sn4_61 sn5_61 11.551961
Rsp4_62 sp4_62 sp5_62 11.551961
Rsn4_62 sn4_62 sn5_62 11.551961
Rsp4_63 sp4_63 sp5_63 11.551961
Rsn4_63 sn4_63 sn5_63 11.551961
Rsp4_64 sp4_64 sp5_64 11.551961
Rsn4_64 sn4_64 sn5_64 11.551961
Rsp4_65 sp4_65 sp5_65 11.551961
Rsn4_65 sn4_65 sn5_65 11.551961
Rsp4_66 sp4_66 sp5_66 11.551961
Rsn4_66 sn4_66 sn5_66 11.551961
Rsp4_67 sp4_67 sp5_67 11.551961
Rsn4_67 sn4_67 sn5_67 11.551961
Rsp4_68 sp4_68 sp5_68 11.551961
Rsn4_68 sn4_68 sn5_68 11.551961
Rsp4_69 sp4_69 sp5_69 11.551961
Rsn4_69 sn4_69 sn5_69 11.551961
Rsp4_70 sp4_70 sp5_70 11.551961
Rsn4_70 sn4_70 sn5_70 11.551961
Rsp4_71 sp4_71 sp5_71 11.551961
Rsn4_71 sn4_71 sn5_71 11.551961
Rsp4_72 sp4_72 sp5_72 11.551961
Rsn4_72 sn4_72 sn5_72 11.551961
Rsp4_73 sp4_73 sp5_73 11.551961
Rsn4_73 sn4_73 sn5_73 11.551961
Rsp4_74 sp4_74 sp5_74 11.551961
Rsn4_74 sn4_74 sn5_74 11.551961
Rsp4_75 sp4_75 sp5_75 11.551961
Rsn4_75 sn4_75 sn5_75 11.551961
Rsp4_76 sp4_76 sp5_76 11.551961
Rsn4_76 sn4_76 sn5_76 11.551961
Rsp4_77 sp4_77 sp5_77 11.551961
Rsn4_77 sn4_77 sn5_77 11.551961
Rsp4_78 sp4_78 sp5_78 11.551961
Rsn4_78 sn4_78 sn5_78 11.551961
Rsp4_79 sp4_79 sp5_79 11.551961
Rsn4_79 sn4_79 sn5_79 11.551961
Rsp4_80 sp4_80 sp5_80 11.551961
Rsn4_80 sn4_80 sn5_80 11.551961
Rsp4_81 sp4_81 sp5_81 11.551961
Rsn4_81 sn4_81 sn5_81 11.551961
Rsp4_82 sp4_82 sp5_82 11.551961
Rsn4_82 sn4_82 sn5_82 11.551961
Rsp4_83 sp4_83 sp5_83 11.551961
Rsn4_83 sn4_83 sn5_83 11.551961
Rsp4_84 sp4_84 sp5_84 11.551961
Rsn4_84 sn4_84 sn5_84 11.551961
Rsp5_1 sp5_1 sp6_1 11.551961
Rsn5_1 sn5_1 sn6_1 11.551961
Rsp5_2 sp5_2 sp6_2 11.551961
Rsn5_2 sn5_2 sn6_2 11.551961
Rsp5_3 sp5_3 sp6_3 11.551961
Rsn5_3 sn5_3 sn6_3 11.551961
Rsp5_4 sp5_4 sp6_4 11.551961
Rsn5_4 sn5_4 sn6_4 11.551961
Rsp5_5 sp5_5 sp6_5 11.551961
Rsn5_5 sn5_5 sn6_5 11.551961
Rsp5_6 sp5_6 sp6_6 11.551961
Rsn5_6 sn5_6 sn6_6 11.551961
Rsp5_7 sp5_7 sp6_7 11.551961
Rsn5_7 sn5_7 sn6_7 11.551961
Rsp5_8 sp5_8 sp6_8 11.551961
Rsn5_8 sn5_8 sn6_8 11.551961
Rsp5_9 sp5_9 sp6_9 11.551961
Rsn5_9 sn5_9 sn6_9 11.551961
Rsp5_10 sp5_10 sp6_10 11.551961
Rsn5_10 sn5_10 sn6_10 11.551961
Rsp5_11 sp5_11 sp6_11 11.551961
Rsn5_11 sn5_11 sn6_11 11.551961
Rsp5_12 sp5_12 sp6_12 11.551961
Rsn5_12 sn5_12 sn6_12 11.551961
Rsp5_13 sp5_13 sp6_13 11.551961
Rsn5_13 sn5_13 sn6_13 11.551961
Rsp5_14 sp5_14 sp6_14 11.551961
Rsn5_14 sn5_14 sn6_14 11.551961
Rsp5_15 sp5_15 sp6_15 11.551961
Rsn5_15 sn5_15 sn6_15 11.551961
Rsp5_16 sp5_16 sp6_16 11.551961
Rsn5_16 sn5_16 sn6_16 11.551961
Rsp5_17 sp5_17 sp6_17 11.551961
Rsn5_17 sn5_17 sn6_17 11.551961
Rsp5_18 sp5_18 sp6_18 11.551961
Rsn5_18 sn5_18 sn6_18 11.551961
Rsp5_19 sp5_19 sp6_19 11.551961
Rsn5_19 sn5_19 sn6_19 11.551961
Rsp5_20 sp5_20 sp6_20 11.551961
Rsn5_20 sn5_20 sn6_20 11.551961
Rsp5_21 sp5_21 sp6_21 11.551961
Rsn5_21 sn5_21 sn6_21 11.551961
Rsp5_22 sp5_22 sp6_22 11.551961
Rsn5_22 sn5_22 sn6_22 11.551961
Rsp5_23 sp5_23 sp6_23 11.551961
Rsn5_23 sn5_23 sn6_23 11.551961
Rsp5_24 sp5_24 sp6_24 11.551961
Rsn5_24 sn5_24 sn6_24 11.551961
Rsp5_25 sp5_25 sp6_25 11.551961
Rsn5_25 sn5_25 sn6_25 11.551961
Rsp5_26 sp5_26 sp6_26 11.551961
Rsn5_26 sn5_26 sn6_26 11.551961
Rsp5_27 sp5_27 sp6_27 11.551961
Rsn5_27 sn5_27 sn6_27 11.551961
Rsp5_28 sp5_28 sp6_28 11.551961
Rsn5_28 sn5_28 sn6_28 11.551961
Rsp5_29 sp5_29 sp6_29 11.551961
Rsn5_29 sn5_29 sn6_29 11.551961
Rsp5_30 sp5_30 sp6_30 11.551961
Rsn5_30 sn5_30 sn6_30 11.551961
Rsp5_31 sp5_31 sp6_31 11.551961
Rsn5_31 sn5_31 sn6_31 11.551961
Rsp5_32 sp5_32 sp6_32 11.551961
Rsn5_32 sn5_32 sn6_32 11.551961
Rsp5_33 sp5_33 sp6_33 11.551961
Rsn5_33 sn5_33 sn6_33 11.551961
Rsp5_34 sp5_34 sp6_34 11.551961
Rsn5_34 sn5_34 sn6_34 11.551961
Rsp5_35 sp5_35 sp6_35 11.551961
Rsn5_35 sn5_35 sn6_35 11.551961
Rsp5_36 sp5_36 sp6_36 11.551961
Rsn5_36 sn5_36 sn6_36 11.551961
Rsp5_37 sp5_37 sp6_37 11.551961
Rsn5_37 sn5_37 sn6_37 11.551961
Rsp5_38 sp5_38 sp6_38 11.551961
Rsn5_38 sn5_38 sn6_38 11.551961
Rsp5_39 sp5_39 sp6_39 11.551961
Rsn5_39 sn5_39 sn6_39 11.551961
Rsp5_40 sp5_40 sp6_40 11.551961
Rsn5_40 sn5_40 sn6_40 11.551961
Rsp5_41 sp5_41 sp6_41 11.551961
Rsn5_41 sn5_41 sn6_41 11.551961
Rsp5_42 sp5_42 sp6_42 11.551961
Rsn5_42 sn5_42 sn6_42 11.551961
Rsp5_43 sp5_43 sp6_43 11.551961
Rsn5_43 sn5_43 sn6_43 11.551961
Rsp5_44 sp5_44 sp6_44 11.551961
Rsn5_44 sn5_44 sn6_44 11.551961
Rsp5_45 sp5_45 sp6_45 11.551961
Rsn5_45 sn5_45 sn6_45 11.551961
Rsp5_46 sp5_46 sp6_46 11.551961
Rsn5_46 sn5_46 sn6_46 11.551961
Rsp5_47 sp5_47 sp6_47 11.551961
Rsn5_47 sn5_47 sn6_47 11.551961
Rsp5_48 sp5_48 sp6_48 11.551961
Rsn5_48 sn5_48 sn6_48 11.551961
Rsp5_49 sp5_49 sp6_49 11.551961
Rsn5_49 sn5_49 sn6_49 11.551961
Rsp5_50 sp5_50 sp6_50 11.551961
Rsn5_50 sn5_50 sn6_50 11.551961
Rsp5_51 sp5_51 sp6_51 11.551961
Rsn5_51 sn5_51 sn6_51 11.551961
Rsp5_52 sp5_52 sp6_52 11.551961
Rsn5_52 sn5_52 sn6_52 11.551961
Rsp5_53 sp5_53 sp6_53 11.551961
Rsn5_53 sn5_53 sn6_53 11.551961
Rsp5_54 sp5_54 sp6_54 11.551961
Rsn5_54 sn5_54 sn6_54 11.551961
Rsp5_55 sp5_55 sp6_55 11.551961
Rsn5_55 sn5_55 sn6_55 11.551961
Rsp5_56 sp5_56 sp6_56 11.551961
Rsn5_56 sn5_56 sn6_56 11.551961
Rsp5_57 sp5_57 sp6_57 11.551961
Rsn5_57 sn5_57 sn6_57 11.551961
Rsp5_58 sp5_58 sp6_58 11.551961
Rsn5_58 sn5_58 sn6_58 11.551961
Rsp5_59 sp5_59 sp6_59 11.551961
Rsn5_59 sn5_59 sn6_59 11.551961
Rsp5_60 sp5_60 sp6_60 11.551961
Rsn5_60 sn5_60 sn6_60 11.551961
Rsp5_61 sp5_61 sp6_61 11.551961
Rsn5_61 sn5_61 sn6_61 11.551961
Rsp5_62 sp5_62 sp6_62 11.551961
Rsn5_62 sn5_62 sn6_62 11.551961
Rsp5_63 sp5_63 sp6_63 11.551961
Rsn5_63 sn5_63 sn6_63 11.551961
Rsp5_64 sp5_64 sp6_64 11.551961
Rsn5_64 sn5_64 sn6_64 11.551961
Rsp5_65 sp5_65 sp6_65 11.551961
Rsn5_65 sn5_65 sn6_65 11.551961
Rsp5_66 sp5_66 sp6_66 11.551961
Rsn5_66 sn5_66 sn6_66 11.551961
Rsp5_67 sp5_67 sp6_67 11.551961
Rsn5_67 sn5_67 sn6_67 11.551961
Rsp5_68 sp5_68 sp6_68 11.551961
Rsn5_68 sn5_68 sn6_68 11.551961
Rsp5_69 sp5_69 sp6_69 11.551961
Rsn5_69 sn5_69 sn6_69 11.551961
Rsp5_70 sp5_70 sp6_70 11.551961
Rsn5_70 sn5_70 sn6_70 11.551961
Rsp5_71 sp5_71 sp6_71 11.551961
Rsn5_71 sn5_71 sn6_71 11.551961
Rsp5_72 sp5_72 sp6_72 11.551961
Rsn5_72 sn5_72 sn6_72 11.551961
Rsp5_73 sp5_73 sp6_73 11.551961
Rsn5_73 sn5_73 sn6_73 11.551961
Rsp5_74 sp5_74 sp6_74 11.551961
Rsn5_74 sn5_74 sn6_74 11.551961
Rsp5_75 sp5_75 sp6_75 11.551961
Rsn5_75 sn5_75 sn6_75 11.551961
Rsp5_76 sp5_76 sp6_76 11.551961
Rsn5_76 sn5_76 sn6_76 11.551961
Rsp5_77 sp5_77 sp6_77 11.551961
Rsn5_77 sn5_77 sn6_77 11.551961
Rsp5_78 sp5_78 sp6_78 11.551961
Rsn5_78 sn5_78 sn6_78 11.551961
Rsp5_79 sp5_79 sp6_79 11.551961
Rsn5_79 sn5_79 sn6_79 11.551961
Rsp5_80 sp5_80 sp6_80 11.551961
Rsn5_80 sn5_80 sn6_80 11.551961
Rsp5_81 sp5_81 sp6_81 11.551961
Rsn5_81 sn5_81 sn6_81 11.551961
Rsp5_82 sp5_82 sp6_82 11.551961
Rsn5_82 sn5_82 sn6_82 11.551961
Rsp5_83 sp5_83 sp6_83 11.551961
Rsn5_83 sn5_83 sn6_83 11.551961
Rsp5_84 sp5_84 sp6_84 11.551961
Rsn5_84 sn5_84 sn6_84 11.551961
Rsp6_1 sp6_1 sp7_1 11.551961
Rsn6_1 sn6_1 sn7_1 11.551961
Rsp6_2 sp6_2 sp7_2 11.551961
Rsn6_2 sn6_2 sn7_2 11.551961
Rsp6_3 sp6_3 sp7_3 11.551961
Rsn6_3 sn6_3 sn7_3 11.551961
Rsp6_4 sp6_4 sp7_4 11.551961
Rsn6_4 sn6_4 sn7_4 11.551961
Rsp6_5 sp6_5 sp7_5 11.551961
Rsn6_5 sn6_5 sn7_5 11.551961
Rsp6_6 sp6_6 sp7_6 11.551961
Rsn6_6 sn6_6 sn7_6 11.551961
Rsp6_7 sp6_7 sp7_7 11.551961
Rsn6_7 sn6_7 sn7_7 11.551961
Rsp6_8 sp6_8 sp7_8 11.551961
Rsn6_8 sn6_8 sn7_8 11.551961
Rsp6_9 sp6_9 sp7_9 11.551961
Rsn6_9 sn6_9 sn7_9 11.551961
Rsp6_10 sp6_10 sp7_10 11.551961
Rsn6_10 sn6_10 sn7_10 11.551961
Rsp6_11 sp6_11 sp7_11 11.551961
Rsn6_11 sn6_11 sn7_11 11.551961
Rsp6_12 sp6_12 sp7_12 11.551961
Rsn6_12 sn6_12 sn7_12 11.551961
Rsp6_13 sp6_13 sp7_13 11.551961
Rsn6_13 sn6_13 sn7_13 11.551961
Rsp6_14 sp6_14 sp7_14 11.551961
Rsn6_14 sn6_14 sn7_14 11.551961
Rsp6_15 sp6_15 sp7_15 11.551961
Rsn6_15 sn6_15 sn7_15 11.551961
Rsp6_16 sp6_16 sp7_16 11.551961
Rsn6_16 sn6_16 sn7_16 11.551961
Rsp6_17 sp6_17 sp7_17 11.551961
Rsn6_17 sn6_17 sn7_17 11.551961
Rsp6_18 sp6_18 sp7_18 11.551961
Rsn6_18 sn6_18 sn7_18 11.551961
Rsp6_19 sp6_19 sp7_19 11.551961
Rsn6_19 sn6_19 sn7_19 11.551961
Rsp6_20 sp6_20 sp7_20 11.551961
Rsn6_20 sn6_20 sn7_20 11.551961
Rsp6_21 sp6_21 sp7_21 11.551961
Rsn6_21 sn6_21 sn7_21 11.551961
Rsp6_22 sp6_22 sp7_22 11.551961
Rsn6_22 sn6_22 sn7_22 11.551961
Rsp6_23 sp6_23 sp7_23 11.551961
Rsn6_23 sn6_23 sn7_23 11.551961
Rsp6_24 sp6_24 sp7_24 11.551961
Rsn6_24 sn6_24 sn7_24 11.551961
Rsp6_25 sp6_25 sp7_25 11.551961
Rsn6_25 sn6_25 sn7_25 11.551961
Rsp6_26 sp6_26 sp7_26 11.551961
Rsn6_26 sn6_26 sn7_26 11.551961
Rsp6_27 sp6_27 sp7_27 11.551961
Rsn6_27 sn6_27 sn7_27 11.551961
Rsp6_28 sp6_28 sp7_28 11.551961
Rsn6_28 sn6_28 sn7_28 11.551961
Rsp6_29 sp6_29 sp7_29 11.551961
Rsn6_29 sn6_29 sn7_29 11.551961
Rsp6_30 sp6_30 sp7_30 11.551961
Rsn6_30 sn6_30 sn7_30 11.551961
Rsp6_31 sp6_31 sp7_31 11.551961
Rsn6_31 sn6_31 sn7_31 11.551961
Rsp6_32 sp6_32 sp7_32 11.551961
Rsn6_32 sn6_32 sn7_32 11.551961
Rsp6_33 sp6_33 sp7_33 11.551961
Rsn6_33 sn6_33 sn7_33 11.551961
Rsp6_34 sp6_34 sp7_34 11.551961
Rsn6_34 sn6_34 sn7_34 11.551961
Rsp6_35 sp6_35 sp7_35 11.551961
Rsn6_35 sn6_35 sn7_35 11.551961
Rsp6_36 sp6_36 sp7_36 11.551961
Rsn6_36 sn6_36 sn7_36 11.551961
Rsp6_37 sp6_37 sp7_37 11.551961
Rsn6_37 sn6_37 sn7_37 11.551961
Rsp6_38 sp6_38 sp7_38 11.551961
Rsn6_38 sn6_38 sn7_38 11.551961
Rsp6_39 sp6_39 sp7_39 11.551961
Rsn6_39 sn6_39 sn7_39 11.551961
Rsp6_40 sp6_40 sp7_40 11.551961
Rsn6_40 sn6_40 sn7_40 11.551961
Rsp6_41 sp6_41 sp7_41 11.551961
Rsn6_41 sn6_41 sn7_41 11.551961
Rsp6_42 sp6_42 sp7_42 11.551961
Rsn6_42 sn6_42 sn7_42 11.551961
Rsp6_43 sp6_43 sp7_43 11.551961
Rsn6_43 sn6_43 sn7_43 11.551961
Rsp6_44 sp6_44 sp7_44 11.551961
Rsn6_44 sn6_44 sn7_44 11.551961
Rsp6_45 sp6_45 sp7_45 11.551961
Rsn6_45 sn6_45 sn7_45 11.551961
Rsp6_46 sp6_46 sp7_46 11.551961
Rsn6_46 sn6_46 sn7_46 11.551961
Rsp6_47 sp6_47 sp7_47 11.551961
Rsn6_47 sn6_47 sn7_47 11.551961
Rsp6_48 sp6_48 sp7_48 11.551961
Rsn6_48 sn6_48 sn7_48 11.551961
Rsp6_49 sp6_49 sp7_49 11.551961
Rsn6_49 sn6_49 sn7_49 11.551961
Rsp6_50 sp6_50 sp7_50 11.551961
Rsn6_50 sn6_50 sn7_50 11.551961
Rsp6_51 sp6_51 sp7_51 11.551961
Rsn6_51 sn6_51 sn7_51 11.551961
Rsp6_52 sp6_52 sp7_52 11.551961
Rsn6_52 sn6_52 sn7_52 11.551961
Rsp6_53 sp6_53 sp7_53 11.551961
Rsn6_53 sn6_53 sn7_53 11.551961
Rsp6_54 sp6_54 sp7_54 11.551961
Rsn6_54 sn6_54 sn7_54 11.551961
Rsp6_55 sp6_55 sp7_55 11.551961
Rsn6_55 sn6_55 sn7_55 11.551961
Rsp6_56 sp6_56 sp7_56 11.551961
Rsn6_56 sn6_56 sn7_56 11.551961
Rsp6_57 sp6_57 sp7_57 11.551961
Rsn6_57 sn6_57 sn7_57 11.551961
Rsp6_58 sp6_58 sp7_58 11.551961
Rsn6_58 sn6_58 sn7_58 11.551961
Rsp6_59 sp6_59 sp7_59 11.551961
Rsn6_59 sn6_59 sn7_59 11.551961
Rsp6_60 sp6_60 sp7_60 11.551961
Rsn6_60 sn6_60 sn7_60 11.551961
Rsp6_61 sp6_61 sp7_61 11.551961
Rsn6_61 sn6_61 sn7_61 11.551961
Rsp6_62 sp6_62 sp7_62 11.551961
Rsn6_62 sn6_62 sn7_62 11.551961
Rsp6_63 sp6_63 sp7_63 11.551961
Rsn6_63 sn6_63 sn7_63 11.551961
Rsp6_64 sp6_64 sp7_64 11.551961
Rsn6_64 sn6_64 sn7_64 11.551961
Rsp6_65 sp6_65 sp7_65 11.551961
Rsn6_65 sn6_65 sn7_65 11.551961
Rsp6_66 sp6_66 sp7_66 11.551961
Rsn6_66 sn6_66 sn7_66 11.551961
Rsp6_67 sp6_67 sp7_67 11.551961
Rsn6_67 sn6_67 sn7_67 11.551961
Rsp6_68 sp6_68 sp7_68 11.551961
Rsn6_68 sn6_68 sn7_68 11.551961
Rsp6_69 sp6_69 sp7_69 11.551961
Rsn6_69 sn6_69 sn7_69 11.551961
Rsp6_70 sp6_70 sp7_70 11.551961
Rsn6_70 sn6_70 sn7_70 11.551961
Rsp6_71 sp6_71 sp7_71 11.551961
Rsn6_71 sn6_71 sn7_71 11.551961
Rsp6_72 sp6_72 sp7_72 11.551961
Rsn6_72 sn6_72 sn7_72 11.551961
Rsp6_73 sp6_73 sp7_73 11.551961
Rsn6_73 sn6_73 sn7_73 11.551961
Rsp6_74 sp6_74 sp7_74 11.551961
Rsn6_74 sn6_74 sn7_74 11.551961
Rsp6_75 sp6_75 sp7_75 11.551961
Rsn6_75 sn6_75 sn7_75 11.551961
Rsp6_76 sp6_76 sp7_76 11.551961
Rsn6_76 sn6_76 sn7_76 11.551961
Rsp6_77 sp6_77 sp7_77 11.551961
Rsn6_77 sn6_77 sn7_77 11.551961
Rsp6_78 sp6_78 sp7_78 11.551961
Rsn6_78 sn6_78 sn7_78 11.551961
Rsp6_79 sp6_79 sp7_79 11.551961
Rsn6_79 sn6_79 sn7_79 11.551961
Rsp6_80 sp6_80 sp7_80 11.551961
Rsn6_80 sn6_80 sn7_80 11.551961
Rsp6_81 sp6_81 sp7_81 11.551961
Rsn6_81 sn6_81 sn7_81 11.551961
Rsp6_82 sp6_82 sp7_82 11.551961
Rsn6_82 sn6_82 sn7_82 11.551961
Rsp6_83 sp6_83 sp7_83 11.551961
Rsn6_83 sn6_83 sn7_83 11.551961
Rsp6_84 sp6_84 sp7_84 11.551961
Rsn6_84 sn6_84 sn7_84 11.551961
Rsp7_1 sp7_1 sp8_1 11.551961
Rsn7_1 sn7_1 sn8_1 11.551961
Rsp7_2 sp7_2 sp8_2 11.551961
Rsn7_2 sn7_2 sn8_2 11.551961
Rsp7_3 sp7_3 sp8_3 11.551961
Rsn7_3 sn7_3 sn8_3 11.551961
Rsp7_4 sp7_4 sp8_4 11.551961
Rsn7_4 sn7_4 sn8_4 11.551961
Rsp7_5 sp7_5 sp8_5 11.551961
Rsn7_5 sn7_5 sn8_5 11.551961
Rsp7_6 sp7_6 sp8_6 11.551961
Rsn7_6 sn7_6 sn8_6 11.551961
Rsp7_7 sp7_7 sp8_7 11.551961
Rsn7_7 sn7_7 sn8_7 11.551961
Rsp7_8 sp7_8 sp8_8 11.551961
Rsn7_8 sn7_8 sn8_8 11.551961
Rsp7_9 sp7_9 sp8_9 11.551961
Rsn7_9 sn7_9 sn8_9 11.551961
Rsp7_10 sp7_10 sp8_10 11.551961
Rsn7_10 sn7_10 sn8_10 11.551961
Rsp7_11 sp7_11 sp8_11 11.551961
Rsn7_11 sn7_11 sn8_11 11.551961
Rsp7_12 sp7_12 sp8_12 11.551961
Rsn7_12 sn7_12 sn8_12 11.551961
Rsp7_13 sp7_13 sp8_13 11.551961
Rsn7_13 sn7_13 sn8_13 11.551961
Rsp7_14 sp7_14 sp8_14 11.551961
Rsn7_14 sn7_14 sn8_14 11.551961
Rsp7_15 sp7_15 sp8_15 11.551961
Rsn7_15 sn7_15 sn8_15 11.551961
Rsp7_16 sp7_16 sp8_16 11.551961
Rsn7_16 sn7_16 sn8_16 11.551961
Rsp7_17 sp7_17 sp8_17 11.551961
Rsn7_17 sn7_17 sn8_17 11.551961
Rsp7_18 sp7_18 sp8_18 11.551961
Rsn7_18 sn7_18 sn8_18 11.551961
Rsp7_19 sp7_19 sp8_19 11.551961
Rsn7_19 sn7_19 sn8_19 11.551961
Rsp7_20 sp7_20 sp8_20 11.551961
Rsn7_20 sn7_20 sn8_20 11.551961
Rsp7_21 sp7_21 sp8_21 11.551961
Rsn7_21 sn7_21 sn8_21 11.551961
Rsp7_22 sp7_22 sp8_22 11.551961
Rsn7_22 sn7_22 sn8_22 11.551961
Rsp7_23 sp7_23 sp8_23 11.551961
Rsn7_23 sn7_23 sn8_23 11.551961
Rsp7_24 sp7_24 sp8_24 11.551961
Rsn7_24 sn7_24 sn8_24 11.551961
Rsp7_25 sp7_25 sp8_25 11.551961
Rsn7_25 sn7_25 sn8_25 11.551961
Rsp7_26 sp7_26 sp8_26 11.551961
Rsn7_26 sn7_26 sn8_26 11.551961
Rsp7_27 sp7_27 sp8_27 11.551961
Rsn7_27 sn7_27 sn8_27 11.551961
Rsp7_28 sp7_28 sp8_28 11.551961
Rsn7_28 sn7_28 sn8_28 11.551961
Rsp7_29 sp7_29 sp8_29 11.551961
Rsn7_29 sn7_29 sn8_29 11.551961
Rsp7_30 sp7_30 sp8_30 11.551961
Rsn7_30 sn7_30 sn8_30 11.551961
Rsp7_31 sp7_31 sp8_31 11.551961
Rsn7_31 sn7_31 sn8_31 11.551961
Rsp7_32 sp7_32 sp8_32 11.551961
Rsn7_32 sn7_32 sn8_32 11.551961
Rsp7_33 sp7_33 sp8_33 11.551961
Rsn7_33 sn7_33 sn8_33 11.551961
Rsp7_34 sp7_34 sp8_34 11.551961
Rsn7_34 sn7_34 sn8_34 11.551961
Rsp7_35 sp7_35 sp8_35 11.551961
Rsn7_35 sn7_35 sn8_35 11.551961
Rsp7_36 sp7_36 sp8_36 11.551961
Rsn7_36 sn7_36 sn8_36 11.551961
Rsp7_37 sp7_37 sp8_37 11.551961
Rsn7_37 sn7_37 sn8_37 11.551961
Rsp7_38 sp7_38 sp8_38 11.551961
Rsn7_38 sn7_38 sn8_38 11.551961
Rsp7_39 sp7_39 sp8_39 11.551961
Rsn7_39 sn7_39 sn8_39 11.551961
Rsp7_40 sp7_40 sp8_40 11.551961
Rsn7_40 sn7_40 sn8_40 11.551961
Rsp7_41 sp7_41 sp8_41 11.551961
Rsn7_41 sn7_41 sn8_41 11.551961
Rsp7_42 sp7_42 sp8_42 11.551961
Rsn7_42 sn7_42 sn8_42 11.551961
Rsp7_43 sp7_43 sp8_43 11.551961
Rsn7_43 sn7_43 sn8_43 11.551961
Rsp7_44 sp7_44 sp8_44 11.551961
Rsn7_44 sn7_44 sn8_44 11.551961
Rsp7_45 sp7_45 sp8_45 11.551961
Rsn7_45 sn7_45 sn8_45 11.551961
Rsp7_46 sp7_46 sp8_46 11.551961
Rsn7_46 sn7_46 sn8_46 11.551961
Rsp7_47 sp7_47 sp8_47 11.551961
Rsn7_47 sn7_47 sn8_47 11.551961
Rsp7_48 sp7_48 sp8_48 11.551961
Rsn7_48 sn7_48 sn8_48 11.551961
Rsp7_49 sp7_49 sp8_49 11.551961
Rsn7_49 sn7_49 sn8_49 11.551961
Rsp7_50 sp7_50 sp8_50 11.551961
Rsn7_50 sn7_50 sn8_50 11.551961
Rsp7_51 sp7_51 sp8_51 11.551961
Rsn7_51 sn7_51 sn8_51 11.551961
Rsp7_52 sp7_52 sp8_52 11.551961
Rsn7_52 sn7_52 sn8_52 11.551961
Rsp7_53 sp7_53 sp8_53 11.551961
Rsn7_53 sn7_53 sn8_53 11.551961
Rsp7_54 sp7_54 sp8_54 11.551961
Rsn7_54 sn7_54 sn8_54 11.551961
Rsp7_55 sp7_55 sp8_55 11.551961
Rsn7_55 sn7_55 sn8_55 11.551961
Rsp7_56 sp7_56 sp8_56 11.551961
Rsn7_56 sn7_56 sn8_56 11.551961
Rsp7_57 sp7_57 sp8_57 11.551961
Rsn7_57 sn7_57 sn8_57 11.551961
Rsp7_58 sp7_58 sp8_58 11.551961
Rsn7_58 sn7_58 sn8_58 11.551961
Rsp7_59 sp7_59 sp8_59 11.551961
Rsn7_59 sn7_59 sn8_59 11.551961
Rsp7_60 sp7_60 sp8_60 11.551961
Rsn7_60 sn7_60 sn8_60 11.551961
Rsp7_61 sp7_61 sp8_61 11.551961
Rsn7_61 sn7_61 sn8_61 11.551961
Rsp7_62 sp7_62 sp8_62 11.551961
Rsn7_62 sn7_62 sn8_62 11.551961
Rsp7_63 sp7_63 sp8_63 11.551961
Rsn7_63 sn7_63 sn8_63 11.551961
Rsp7_64 sp7_64 sp8_64 11.551961
Rsn7_64 sn7_64 sn8_64 11.551961
Rsp7_65 sp7_65 sp8_65 11.551961
Rsn7_65 sn7_65 sn8_65 11.551961
Rsp7_66 sp7_66 sp8_66 11.551961
Rsn7_66 sn7_66 sn8_66 11.551961
Rsp7_67 sp7_67 sp8_67 11.551961
Rsn7_67 sn7_67 sn8_67 11.551961
Rsp7_68 sp7_68 sp8_68 11.551961
Rsn7_68 sn7_68 sn8_68 11.551961
Rsp7_69 sp7_69 sp8_69 11.551961
Rsn7_69 sn7_69 sn8_69 11.551961
Rsp7_70 sp7_70 sp8_70 11.551961
Rsn7_70 sn7_70 sn8_70 11.551961
Rsp7_71 sp7_71 sp8_71 11.551961
Rsn7_71 sn7_71 sn8_71 11.551961
Rsp7_72 sp7_72 sp8_72 11.551961
Rsn7_72 sn7_72 sn8_72 11.551961
Rsp7_73 sp7_73 sp8_73 11.551961
Rsn7_73 sn7_73 sn8_73 11.551961
Rsp7_74 sp7_74 sp8_74 11.551961
Rsn7_74 sn7_74 sn8_74 11.551961
Rsp7_75 sp7_75 sp8_75 11.551961
Rsn7_75 sn7_75 sn8_75 11.551961
Rsp7_76 sp7_76 sp8_76 11.551961
Rsn7_76 sn7_76 sn8_76 11.551961
Rsp7_77 sp7_77 sp8_77 11.551961
Rsn7_77 sn7_77 sn8_77 11.551961
Rsp7_78 sp7_78 sp8_78 11.551961
Rsn7_78 sn7_78 sn8_78 11.551961
Rsp7_79 sp7_79 sp8_79 11.551961
Rsn7_79 sn7_79 sn8_79 11.551961
Rsp7_80 sp7_80 sp8_80 11.551961
Rsn7_80 sn7_80 sn8_80 11.551961
Rsp7_81 sp7_81 sp8_81 11.551961
Rsn7_81 sn7_81 sn8_81 11.551961
Rsp7_82 sp7_82 sp8_82 11.551961
Rsn7_82 sn7_82 sn8_82 11.551961
Rsp7_83 sp7_83 sp8_83 11.551961
Rsn7_83 sn7_83 sn8_83 11.551961
Rsp7_84 sp7_84 sp8_84 11.551961
Rsn7_84 sn7_84 sn8_84 11.551961
Rsp8_1 sp8_1 sp9_1 11.551961
Rsn8_1 sn8_1 sn9_1 11.551961
Rsp8_2 sp8_2 sp9_2 11.551961
Rsn8_2 sn8_2 sn9_2 11.551961
Rsp8_3 sp8_3 sp9_3 11.551961
Rsn8_3 sn8_3 sn9_3 11.551961
Rsp8_4 sp8_4 sp9_4 11.551961
Rsn8_4 sn8_4 sn9_4 11.551961
Rsp8_5 sp8_5 sp9_5 11.551961
Rsn8_5 sn8_5 sn9_5 11.551961
Rsp8_6 sp8_6 sp9_6 11.551961
Rsn8_6 sn8_6 sn9_6 11.551961
Rsp8_7 sp8_7 sp9_7 11.551961
Rsn8_7 sn8_7 sn9_7 11.551961
Rsp8_8 sp8_8 sp9_8 11.551961
Rsn8_8 sn8_8 sn9_8 11.551961
Rsp8_9 sp8_9 sp9_9 11.551961
Rsn8_9 sn8_9 sn9_9 11.551961
Rsp8_10 sp8_10 sp9_10 11.551961
Rsn8_10 sn8_10 sn9_10 11.551961
Rsp8_11 sp8_11 sp9_11 11.551961
Rsn8_11 sn8_11 sn9_11 11.551961
Rsp8_12 sp8_12 sp9_12 11.551961
Rsn8_12 sn8_12 sn9_12 11.551961
Rsp8_13 sp8_13 sp9_13 11.551961
Rsn8_13 sn8_13 sn9_13 11.551961
Rsp8_14 sp8_14 sp9_14 11.551961
Rsn8_14 sn8_14 sn9_14 11.551961
Rsp8_15 sp8_15 sp9_15 11.551961
Rsn8_15 sn8_15 sn9_15 11.551961
Rsp8_16 sp8_16 sp9_16 11.551961
Rsn8_16 sn8_16 sn9_16 11.551961
Rsp8_17 sp8_17 sp9_17 11.551961
Rsn8_17 sn8_17 sn9_17 11.551961
Rsp8_18 sp8_18 sp9_18 11.551961
Rsn8_18 sn8_18 sn9_18 11.551961
Rsp8_19 sp8_19 sp9_19 11.551961
Rsn8_19 sn8_19 sn9_19 11.551961
Rsp8_20 sp8_20 sp9_20 11.551961
Rsn8_20 sn8_20 sn9_20 11.551961
Rsp8_21 sp8_21 sp9_21 11.551961
Rsn8_21 sn8_21 sn9_21 11.551961
Rsp8_22 sp8_22 sp9_22 11.551961
Rsn8_22 sn8_22 sn9_22 11.551961
Rsp8_23 sp8_23 sp9_23 11.551961
Rsn8_23 sn8_23 sn9_23 11.551961
Rsp8_24 sp8_24 sp9_24 11.551961
Rsn8_24 sn8_24 sn9_24 11.551961
Rsp8_25 sp8_25 sp9_25 11.551961
Rsn8_25 sn8_25 sn9_25 11.551961
Rsp8_26 sp8_26 sp9_26 11.551961
Rsn8_26 sn8_26 sn9_26 11.551961
Rsp8_27 sp8_27 sp9_27 11.551961
Rsn8_27 sn8_27 sn9_27 11.551961
Rsp8_28 sp8_28 sp9_28 11.551961
Rsn8_28 sn8_28 sn9_28 11.551961
Rsp8_29 sp8_29 sp9_29 11.551961
Rsn8_29 sn8_29 sn9_29 11.551961
Rsp8_30 sp8_30 sp9_30 11.551961
Rsn8_30 sn8_30 sn9_30 11.551961
Rsp8_31 sp8_31 sp9_31 11.551961
Rsn8_31 sn8_31 sn9_31 11.551961
Rsp8_32 sp8_32 sp9_32 11.551961
Rsn8_32 sn8_32 sn9_32 11.551961
Rsp8_33 sp8_33 sp9_33 11.551961
Rsn8_33 sn8_33 sn9_33 11.551961
Rsp8_34 sp8_34 sp9_34 11.551961
Rsn8_34 sn8_34 sn9_34 11.551961
Rsp8_35 sp8_35 sp9_35 11.551961
Rsn8_35 sn8_35 sn9_35 11.551961
Rsp8_36 sp8_36 sp9_36 11.551961
Rsn8_36 sn8_36 sn9_36 11.551961
Rsp8_37 sp8_37 sp9_37 11.551961
Rsn8_37 sn8_37 sn9_37 11.551961
Rsp8_38 sp8_38 sp9_38 11.551961
Rsn8_38 sn8_38 sn9_38 11.551961
Rsp8_39 sp8_39 sp9_39 11.551961
Rsn8_39 sn8_39 sn9_39 11.551961
Rsp8_40 sp8_40 sp9_40 11.551961
Rsn8_40 sn8_40 sn9_40 11.551961
Rsp8_41 sp8_41 sp9_41 11.551961
Rsn8_41 sn8_41 sn9_41 11.551961
Rsp8_42 sp8_42 sp9_42 11.551961
Rsn8_42 sn8_42 sn9_42 11.551961
Rsp8_43 sp8_43 sp9_43 11.551961
Rsn8_43 sn8_43 sn9_43 11.551961
Rsp8_44 sp8_44 sp9_44 11.551961
Rsn8_44 sn8_44 sn9_44 11.551961
Rsp8_45 sp8_45 sp9_45 11.551961
Rsn8_45 sn8_45 sn9_45 11.551961
Rsp8_46 sp8_46 sp9_46 11.551961
Rsn8_46 sn8_46 sn9_46 11.551961
Rsp8_47 sp8_47 sp9_47 11.551961
Rsn8_47 sn8_47 sn9_47 11.551961
Rsp8_48 sp8_48 sp9_48 11.551961
Rsn8_48 sn8_48 sn9_48 11.551961
Rsp8_49 sp8_49 sp9_49 11.551961
Rsn8_49 sn8_49 sn9_49 11.551961
Rsp8_50 sp8_50 sp9_50 11.551961
Rsn8_50 sn8_50 sn9_50 11.551961
Rsp8_51 sp8_51 sp9_51 11.551961
Rsn8_51 sn8_51 sn9_51 11.551961
Rsp8_52 sp8_52 sp9_52 11.551961
Rsn8_52 sn8_52 sn9_52 11.551961
Rsp8_53 sp8_53 sp9_53 11.551961
Rsn8_53 sn8_53 sn9_53 11.551961
Rsp8_54 sp8_54 sp9_54 11.551961
Rsn8_54 sn8_54 sn9_54 11.551961
Rsp8_55 sp8_55 sp9_55 11.551961
Rsn8_55 sn8_55 sn9_55 11.551961
Rsp8_56 sp8_56 sp9_56 11.551961
Rsn8_56 sn8_56 sn9_56 11.551961
Rsp8_57 sp8_57 sp9_57 11.551961
Rsn8_57 sn8_57 sn9_57 11.551961
Rsp8_58 sp8_58 sp9_58 11.551961
Rsn8_58 sn8_58 sn9_58 11.551961
Rsp8_59 sp8_59 sp9_59 11.551961
Rsn8_59 sn8_59 sn9_59 11.551961
Rsp8_60 sp8_60 sp9_60 11.551961
Rsn8_60 sn8_60 sn9_60 11.551961
Rsp8_61 sp8_61 sp9_61 11.551961
Rsn8_61 sn8_61 sn9_61 11.551961
Rsp8_62 sp8_62 sp9_62 11.551961
Rsn8_62 sn8_62 sn9_62 11.551961
Rsp8_63 sp8_63 sp9_63 11.551961
Rsn8_63 sn8_63 sn9_63 11.551961
Rsp8_64 sp8_64 sp9_64 11.551961
Rsn8_64 sn8_64 sn9_64 11.551961
Rsp8_65 sp8_65 sp9_65 11.551961
Rsn8_65 sn8_65 sn9_65 11.551961
Rsp8_66 sp8_66 sp9_66 11.551961
Rsn8_66 sn8_66 sn9_66 11.551961
Rsp8_67 sp8_67 sp9_67 11.551961
Rsn8_67 sn8_67 sn9_67 11.551961
Rsp8_68 sp8_68 sp9_68 11.551961
Rsn8_68 sn8_68 sn9_68 11.551961
Rsp8_69 sp8_69 sp9_69 11.551961
Rsn8_69 sn8_69 sn9_69 11.551961
Rsp8_70 sp8_70 sp9_70 11.551961
Rsn8_70 sn8_70 sn9_70 11.551961
Rsp8_71 sp8_71 sp9_71 11.551961
Rsn8_71 sn8_71 sn9_71 11.551961
Rsp8_72 sp8_72 sp9_72 11.551961
Rsn8_72 sn8_72 sn9_72 11.551961
Rsp8_73 sp8_73 sp9_73 11.551961
Rsn8_73 sn8_73 sn9_73 11.551961
Rsp8_74 sp8_74 sp9_74 11.551961
Rsn8_74 sn8_74 sn9_74 11.551961
Rsp8_75 sp8_75 sp9_75 11.551961
Rsn8_75 sn8_75 sn9_75 11.551961
Rsp8_76 sp8_76 sp9_76 11.551961
Rsn8_76 sn8_76 sn9_76 11.551961
Rsp8_77 sp8_77 sp9_77 11.551961
Rsn8_77 sn8_77 sn9_77 11.551961
Rsp8_78 sp8_78 sp9_78 11.551961
Rsn8_78 sn8_78 sn9_78 11.551961
Rsp8_79 sp8_79 sp9_79 11.551961
Rsn8_79 sn8_79 sn9_79 11.551961
Rsp8_80 sp8_80 sp9_80 11.551961
Rsn8_80 sn8_80 sn9_80 11.551961
Rsp8_81 sp8_81 sp9_81 11.551961
Rsn8_81 sn8_81 sn9_81 11.551961
Rsp8_82 sp8_82 sp9_82 11.551961
Rsn8_82 sn8_82 sn9_82 11.551961
Rsp8_83 sp8_83 sp9_83 11.551961
Rsn8_83 sn8_83 sn9_83 11.551961
Rsp8_84 sp8_84 sp9_84 11.551961
Rsn8_84 sn8_84 sn9_84 11.551961
Rsp9_1 sp9_1 sp10_1 11.551961
Rsn9_1 sn9_1 sn10_1 11.551961
Rsp9_2 sp9_2 sp10_2 11.551961
Rsn9_2 sn9_2 sn10_2 11.551961
Rsp9_3 sp9_3 sp10_3 11.551961
Rsn9_3 sn9_3 sn10_3 11.551961
Rsp9_4 sp9_4 sp10_4 11.551961
Rsn9_4 sn9_4 sn10_4 11.551961
Rsp9_5 sp9_5 sp10_5 11.551961
Rsn9_5 sn9_5 sn10_5 11.551961
Rsp9_6 sp9_6 sp10_6 11.551961
Rsn9_6 sn9_6 sn10_6 11.551961
Rsp9_7 sp9_7 sp10_7 11.551961
Rsn9_7 sn9_7 sn10_7 11.551961
Rsp9_8 sp9_8 sp10_8 11.551961
Rsn9_8 sn9_8 sn10_8 11.551961
Rsp9_9 sp9_9 sp10_9 11.551961
Rsn9_9 sn9_9 sn10_9 11.551961
Rsp9_10 sp9_10 sp10_10 11.551961
Rsn9_10 sn9_10 sn10_10 11.551961
Rsp9_11 sp9_11 sp10_11 11.551961
Rsn9_11 sn9_11 sn10_11 11.551961
Rsp9_12 sp9_12 sp10_12 11.551961
Rsn9_12 sn9_12 sn10_12 11.551961
Rsp9_13 sp9_13 sp10_13 11.551961
Rsn9_13 sn9_13 sn10_13 11.551961
Rsp9_14 sp9_14 sp10_14 11.551961
Rsn9_14 sn9_14 sn10_14 11.551961
Rsp9_15 sp9_15 sp10_15 11.551961
Rsn9_15 sn9_15 sn10_15 11.551961
Rsp9_16 sp9_16 sp10_16 11.551961
Rsn9_16 sn9_16 sn10_16 11.551961
Rsp9_17 sp9_17 sp10_17 11.551961
Rsn9_17 sn9_17 sn10_17 11.551961
Rsp9_18 sp9_18 sp10_18 11.551961
Rsn9_18 sn9_18 sn10_18 11.551961
Rsp9_19 sp9_19 sp10_19 11.551961
Rsn9_19 sn9_19 sn10_19 11.551961
Rsp9_20 sp9_20 sp10_20 11.551961
Rsn9_20 sn9_20 sn10_20 11.551961
Rsp9_21 sp9_21 sp10_21 11.551961
Rsn9_21 sn9_21 sn10_21 11.551961
Rsp9_22 sp9_22 sp10_22 11.551961
Rsn9_22 sn9_22 sn10_22 11.551961
Rsp9_23 sp9_23 sp10_23 11.551961
Rsn9_23 sn9_23 sn10_23 11.551961
Rsp9_24 sp9_24 sp10_24 11.551961
Rsn9_24 sn9_24 sn10_24 11.551961
Rsp9_25 sp9_25 sp10_25 11.551961
Rsn9_25 sn9_25 sn10_25 11.551961
Rsp9_26 sp9_26 sp10_26 11.551961
Rsn9_26 sn9_26 sn10_26 11.551961
Rsp9_27 sp9_27 sp10_27 11.551961
Rsn9_27 sn9_27 sn10_27 11.551961
Rsp9_28 sp9_28 sp10_28 11.551961
Rsn9_28 sn9_28 sn10_28 11.551961
Rsp9_29 sp9_29 sp10_29 11.551961
Rsn9_29 sn9_29 sn10_29 11.551961
Rsp9_30 sp9_30 sp10_30 11.551961
Rsn9_30 sn9_30 sn10_30 11.551961
Rsp9_31 sp9_31 sp10_31 11.551961
Rsn9_31 sn9_31 sn10_31 11.551961
Rsp9_32 sp9_32 sp10_32 11.551961
Rsn9_32 sn9_32 sn10_32 11.551961
Rsp9_33 sp9_33 sp10_33 11.551961
Rsn9_33 sn9_33 sn10_33 11.551961
Rsp9_34 sp9_34 sp10_34 11.551961
Rsn9_34 sn9_34 sn10_34 11.551961
Rsp9_35 sp9_35 sp10_35 11.551961
Rsn9_35 sn9_35 sn10_35 11.551961
Rsp9_36 sp9_36 sp10_36 11.551961
Rsn9_36 sn9_36 sn10_36 11.551961
Rsp9_37 sp9_37 sp10_37 11.551961
Rsn9_37 sn9_37 sn10_37 11.551961
Rsp9_38 sp9_38 sp10_38 11.551961
Rsn9_38 sn9_38 sn10_38 11.551961
Rsp9_39 sp9_39 sp10_39 11.551961
Rsn9_39 sn9_39 sn10_39 11.551961
Rsp9_40 sp9_40 sp10_40 11.551961
Rsn9_40 sn9_40 sn10_40 11.551961
Rsp9_41 sp9_41 sp10_41 11.551961
Rsn9_41 sn9_41 sn10_41 11.551961
Rsp9_42 sp9_42 sp10_42 11.551961
Rsn9_42 sn9_42 sn10_42 11.551961
Rsp9_43 sp9_43 sp10_43 11.551961
Rsn9_43 sn9_43 sn10_43 11.551961
Rsp9_44 sp9_44 sp10_44 11.551961
Rsn9_44 sn9_44 sn10_44 11.551961
Rsp9_45 sp9_45 sp10_45 11.551961
Rsn9_45 sn9_45 sn10_45 11.551961
Rsp9_46 sp9_46 sp10_46 11.551961
Rsn9_46 sn9_46 sn10_46 11.551961
Rsp9_47 sp9_47 sp10_47 11.551961
Rsn9_47 sn9_47 sn10_47 11.551961
Rsp9_48 sp9_48 sp10_48 11.551961
Rsn9_48 sn9_48 sn10_48 11.551961
Rsp9_49 sp9_49 sp10_49 11.551961
Rsn9_49 sn9_49 sn10_49 11.551961
Rsp9_50 sp9_50 sp10_50 11.551961
Rsn9_50 sn9_50 sn10_50 11.551961
Rsp9_51 sp9_51 sp10_51 11.551961
Rsn9_51 sn9_51 sn10_51 11.551961
Rsp9_52 sp9_52 sp10_52 11.551961
Rsn9_52 sn9_52 sn10_52 11.551961
Rsp9_53 sp9_53 sp10_53 11.551961
Rsn9_53 sn9_53 sn10_53 11.551961
Rsp9_54 sp9_54 sp10_54 11.551961
Rsn9_54 sn9_54 sn10_54 11.551961
Rsp9_55 sp9_55 sp10_55 11.551961
Rsn9_55 sn9_55 sn10_55 11.551961
Rsp9_56 sp9_56 sp10_56 11.551961
Rsn9_56 sn9_56 sn10_56 11.551961
Rsp9_57 sp9_57 sp10_57 11.551961
Rsn9_57 sn9_57 sn10_57 11.551961
Rsp9_58 sp9_58 sp10_58 11.551961
Rsn9_58 sn9_58 sn10_58 11.551961
Rsp9_59 sp9_59 sp10_59 11.551961
Rsn9_59 sn9_59 sn10_59 11.551961
Rsp9_60 sp9_60 sp10_60 11.551961
Rsn9_60 sn9_60 sn10_60 11.551961
Rsp9_61 sp9_61 sp10_61 11.551961
Rsn9_61 sn9_61 sn10_61 11.551961
Rsp9_62 sp9_62 sp10_62 11.551961
Rsn9_62 sn9_62 sn10_62 11.551961
Rsp9_63 sp9_63 sp10_63 11.551961
Rsn9_63 sn9_63 sn10_63 11.551961
Rsp9_64 sp9_64 sp10_64 11.551961
Rsn9_64 sn9_64 sn10_64 11.551961
Rsp9_65 sp9_65 sp10_65 11.551961
Rsn9_65 sn9_65 sn10_65 11.551961
Rsp9_66 sp9_66 sp10_66 11.551961
Rsn9_66 sn9_66 sn10_66 11.551961
Rsp9_67 sp9_67 sp10_67 11.551961
Rsn9_67 sn9_67 sn10_67 11.551961
Rsp9_68 sp9_68 sp10_68 11.551961
Rsn9_68 sn9_68 sn10_68 11.551961
Rsp9_69 sp9_69 sp10_69 11.551961
Rsn9_69 sn9_69 sn10_69 11.551961
Rsp9_70 sp9_70 sp10_70 11.551961
Rsn9_70 sn9_70 sn10_70 11.551961
Rsp9_71 sp9_71 sp10_71 11.551961
Rsn9_71 sn9_71 sn10_71 11.551961
Rsp9_72 sp9_72 sp10_72 11.551961
Rsn9_72 sn9_72 sn10_72 11.551961
Rsp9_73 sp9_73 sp10_73 11.551961
Rsn9_73 sn9_73 sn10_73 11.551961
Rsp9_74 sp9_74 sp10_74 11.551961
Rsn9_74 sn9_74 sn10_74 11.551961
Rsp9_75 sp9_75 sp10_75 11.551961
Rsn9_75 sn9_75 sn10_75 11.551961
Rsp9_76 sp9_76 sp10_76 11.551961
Rsn9_76 sn9_76 sn10_76 11.551961
Rsp9_77 sp9_77 sp10_77 11.551961
Rsn9_77 sn9_77 sn10_77 11.551961
Rsp9_78 sp9_78 sp10_78 11.551961
Rsn9_78 sn9_78 sn10_78 11.551961
Rsp9_79 sp9_79 sp10_79 11.551961
Rsn9_79 sn9_79 sn10_79 11.551961
Rsp9_80 sp9_80 sp10_80 11.551961
Rsn9_80 sn9_80 sn10_80 11.551961
Rsp9_81 sp9_81 sp10_81 11.551961
Rsn9_81 sn9_81 sn10_81 11.551961
Rsp9_82 sp9_82 sp10_82 11.551961
Rsn9_82 sn9_82 sn10_82 11.551961
Rsp9_83 sp9_83 sp10_83 11.551961
Rsn9_83 sn9_83 sn10_83 11.551961
Rsp9_84 sp9_84 sp10_84 11.551961
Rsn9_84 sn9_84 sn10_84 11.551961
Rsp10_1 sp10_1 sp11_1 11.551961
Rsn10_1 sn10_1 sn11_1 11.551961
Rsp10_2 sp10_2 sp11_2 11.551961
Rsn10_2 sn10_2 sn11_2 11.551961
Rsp10_3 sp10_3 sp11_3 11.551961
Rsn10_3 sn10_3 sn11_3 11.551961
Rsp10_4 sp10_4 sp11_4 11.551961
Rsn10_4 sn10_4 sn11_4 11.551961
Rsp10_5 sp10_5 sp11_5 11.551961
Rsn10_5 sn10_5 sn11_5 11.551961
Rsp10_6 sp10_6 sp11_6 11.551961
Rsn10_6 sn10_6 sn11_6 11.551961
Rsp10_7 sp10_7 sp11_7 11.551961
Rsn10_7 sn10_7 sn11_7 11.551961
Rsp10_8 sp10_8 sp11_8 11.551961
Rsn10_8 sn10_8 sn11_8 11.551961
Rsp10_9 sp10_9 sp11_9 11.551961
Rsn10_9 sn10_9 sn11_9 11.551961
Rsp10_10 sp10_10 sp11_10 11.551961
Rsn10_10 sn10_10 sn11_10 11.551961
Rsp10_11 sp10_11 sp11_11 11.551961
Rsn10_11 sn10_11 sn11_11 11.551961
Rsp10_12 sp10_12 sp11_12 11.551961
Rsn10_12 sn10_12 sn11_12 11.551961
Rsp10_13 sp10_13 sp11_13 11.551961
Rsn10_13 sn10_13 sn11_13 11.551961
Rsp10_14 sp10_14 sp11_14 11.551961
Rsn10_14 sn10_14 sn11_14 11.551961
Rsp10_15 sp10_15 sp11_15 11.551961
Rsn10_15 sn10_15 sn11_15 11.551961
Rsp10_16 sp10_16 sp11_16 11.551961
Rsn10_16 sn10_16 sn11_16 11.551961
Rsp10_17 sp10_17 sp11_17 11.551961
Rsn10_17 sn10_17 sn11_17 11.551961
Rsp10_18 sp10_18 sp11_18 11.551961
Rsn10_18 sn10_18 sn11_18 11.551961
Rsp10_19 sp10_19 sp11_19 11.551961
Rsn10_19 sn10_19 sn11_19 11.551961
Rsp10_20 sp10_20 sp11_20 11.551961
Rsn10_20 sn10_20 sn11_20 11.551961
Rsp10_21 sp10_21 sp11_21 11.551961
Rsn10_21 sn10_21 sn11_21 11.551961
Rsp10_22 sp10_22 sp11_22 11.551961
Rsn10_22 sn10_22 sn11_22 11.551961
Rsp10_23 sp10_23 sp11_23 11.551961
Rsn10_23 sn10_23 sn11_23 11.551961
Rsp10_24 sp10_24 sp11_24 11.551961
Rsn10_24 sn10_24 sn11_24 11.551961
Rsp10_25 sp10_25 sp11_25 11.551961
Rsn10_25 sn10_25 sn11_25 11.551961
Rsp10_26 sp10_26 sp11_26 11.551961
Rsn10_26 sn10_26 sn11_26 11.551961
Rsp10_27 sp10_27 sp11_27 11.551961
Rsn10_27 sn10_27 sn11_27 11.551961
Rsp10_28 sp10_28 sp11_28 11.551961
Rsn10_28 sn10_28 sn11_28 11.551961
Rsp10_29 sp10_29 sp11_29 11.551961
Rsn10_29 sn10_29 sn11_29 11.551961
Rsp10_30 sp10_30 sp11_30 11.551961
Rsn10_30 sn10_30 sn11_30 11.551961
Rsp10_31 sp10_31 sp11_31 11.551961
Rsn10_31 sn10_31 sn11_31 11.551961
Rsp10_32 sp10_32 sp11_32 11.551961
Rsn10_32 sn10_32 sn11_32 11.551961
Rsp10_33 sp10_33 sp11_33 11.551961
Rsn10_33 sn10_33 sn11_33 11.551961
Rsp10_34 sp10_34 sp11_34 11.551961
Rsn10_34 sn10_34 sn11_34 11.551961
Rsp10_35 sp10_35 sp11_35 11.551961
Rsn10_35 sn10_35 sn11_35 11.551961
Rsp10_36 sp10_36 sp11_36 11.551961
Rsn10_36 sn10_36 sn11_36 11.551961
Rsp10_37 sp10_37 sp11_37 11.551961
Rsn10_37 sn10_37 sn11_37 11.551961
Rsp10_38 sp10_38 sp11_38 11.551961
Rsn10_38 sn10_38 sn11_38 11.551961
Rsp10_39 sp10_39 sp11_39 11.551961
Rsn10_39 sn10_39 sn11_39 11.551961
Rsp10_40 sp10_40 sp11_40 11.551961
Rsn10_40 sn10_40 sn11_40 11.551961
Rsp10_41 sp10_41 sp11_41 11.551961
Rsn10_41 sn10_41 sn11_41 11.551961
Rsp10_42 sp10_42 sp11_42 11.551961
Rsn10_42 sn10_42 sn11_42 11.551961
Rsp10_43 sp10_43 sp11_43 11.551961
Rsn10_43 sn10_43 sn11_43 11.551961
Rsp10_44 sp10_44 sp11_44 11.551961
Rsn10_44 sn10_44 sn11_44 11.551961
Rsp10_45 sp10_45 sp11_45 11.551961
Rsn10_45 sn10_45 sn11_45 11.551961
Rsp10_46 sp10_46 sp11_46 11.551961
Rsn10_46 sn10_46 sn11_46 11.551961
Rsp10_47 sp10_47 sp11_47 11.551961
Rsn10_47 sn10_47 sn11_47 11.551961
Rsp10_48 sp10_48 sp11_48 11.551961
Rsn10_48 sn10_48 sn11_48 11.551961
Rsp10_49 sp10_49 sp11_49 11.551961
Rsn10_49 sn10_49 sn11_49 11.551961
Rsp10_50 sp10_50 sp11_50 11.551961
Rsn10_50 sn10_50 sn11_50 11.551961
Rsp10_51 sp10_51 sp11_51 11.551961
Rsn10_51 sn10_51 sn11_51 11.551961
Rsp10_52 sp10_52 sp11_52 11.551961
Rsn10_52 sn10_52 sn11_52 11.551961
Rsp10_53 sp10_53 sp11_53 11.551961
Rsn10_53 sn10_53 sn11_53 11.551961
Rsp10_54 sp10_54 sp11_54 11.551961
Rsn10_54 sn10_54 sn11_54 11.551961
Rsp10_55 sp10_55 sp11_55 11.551961
Rsn10_55 sn10_55 sn11_55 11.551961
Rsp10_56 sp10_56 sp11_56 11.551961
Rsn10_56 sn10_56 sn11_56 11.551961
Rsp10_57 sp10_57 sp11_57 11.551961
Rsn10_57 sn10_57 sn11_57 11.551961
Rsp10_58 sp10_58 sp11_58 11.551961
Rsn10_58 sn10_58 sn11_58 11.551961
Rsp10_59 sp10_59 sp11_59 11.551961
Rsn10_59 sn10_59 sn11_59 11.551961
Rsp10_60 sp10_60 sp11_60 11.551961
Rsn10_60 sn10_60 sn11_60 11.551961
Rsp10_61 sp10_61 sp11_61 11.551961
Rsn10_61 sn10_61 sn11_61 11.551961
Rsp10_62 sp10_62 sp11_62 11.551961
Rsn10_62 sn10_62 sn11_62 11.551961
Rsp10_63 sp10_63 sp11_63 11.551961
Rsn10_63 sn10_63 sn11_63 11.551961
Rsp10_64 sp10_64 sp11_64 11.551961
Rsn10_64 sn10_64 sn11_64 11.551961
Rsp10_65 sp10_65 sp11_65 11.551961
Rsn10_65 sn10_65 sn11_65 11.551961
Rsp10_66 sp10_66 sp11_66 11.551961
Rsn10_66 sn10_66 sn11_66 11.551961
Rsp10_67 sp10_67 sp11_67 11.551961
Rsn10_67 sn10_67 sn11_67 11.551961
Rsp10_68 sp10_68 sp11_68 11.551961
Rsn10_68 sn10_68 sn11_68 11.551961
Rsp10_69 sp10_69 sp11_69 11.551961
Rsn10_69 sn10_69 sn11_69 11.551961
Rsp10_70 sp10_70 sp11_70 11.551961
Rsn10_70 sn10_70 sn11_70 11.551961
Rsp10_71 sp10_71 sp11_71 11.551961
Rsn10_71 sn10_71 sn11_71 11.551961
Rsp10_72 sp10_72 sp11_72 11.551961
Rsn10_72 sn10_72 sn11_72 11.551961
Rsp10_73 sp10_73 sp11_73 11.551961
Rsn10_73 sn10_73 sn11_73 11.551961
Rsp10_74 sp10_74 sp11_74 11.551961
Rsn10_74 sn10_74 sn11_74 11.551961
Rsp10_75 sp10_75 sp11_75 11.551961
Rsn10_75 sn10_75 sn11_75 11.551961
Rsp10_76 sp10_76 sp11_76 11.551961
Rsn10_76 sn10_76 sn11_76 11.551961
Rsp10_77 sp10_77 sp11_77 11.551961
Rsn10_77 sn10_77 sn11_77 11.551961
Rsp10_78 sp10_78 sp11_78 11.551961
Rsn10_78 sn10_78 sn11_78 11.551961
Rsp10_79 sp10_79 sp11_79 11.551961
Rsn10_79 sn10_79 sn11_79 11.551961
Rsp10_80 sp10_80 sp11_80 11.551961
Rsn10_80 sn10_80 sn11_80 11.551961
Rsp10_81 sp10_81 sp11_81 11.551961
Rsn10_81 sn10_81 sn11_81 11.551961
Rsp10_82 sp10_82 sp11_82 11.551961
Rsn10_82 sn10_82 sn11_82 11.551961
Rsp10_83 sp10_83 sp11_83 11.551961
Rsn10_83 sn10_83 sn11_83 11.551961
Rsp10_84 sp10_84 sp11_84 11.551961
Rsn10_84 sn10_84 sn11_84 11.551961
Rsp11_1 sp11_1 sp12_1 11.551961
Rsn11_1 sn11_1 sn12_1 11.551961
Rsp11_2 sp11_2 sp12_2 11.551961
Rsn11_2 sn11_2 sn12_2 11.551961
Rsp11_3 sp11_3 sp12_3 11.551961
Rsn11_3 sn11_3 sn12_3 11.551961
Rsp11_4 sp11_4 sp12_4 11.551961
Rsn11_4 sn11_4 sn12_4 11.551961
Rsp11_5 sp11_5 sp12_5 11.551961
Rsn11_5 sn11_5 sn12_5 11.551961
Rsp11_6 sp11_6 sp12_6 11.551961
Rsn11_6 sn11_6 sn12_6 11.551961
Rsp11_7 sp11_7 sp12_7 11.551961
Rsn11_7 sn11_7 sn12_7 11.551961
Rsp11_8 sp11_8 sp12_8 11.551961
Rsn11_8 sn11_8 sn12_8 11.551961
Rsp11_9 sp11_9 sp12_9 11.551961
Rsn11_9 sn11_9 sn12_9 11.551961
Rsp11_10 sp11_10 sp12_10 11.551961
Rsn11_10 sn11_10 sn12_10 11.551961
Rsp11_11 sp11_11 sp12_11 11.551961
Rsn11_11 sn11_11 sn12_11 11.551961
Rsp11_12 sp11_12 sp12_12 11.551961
Rsn11_12 sn11_12 sn12_12 11.551961
Rsp11_13 sp11_13 sp12_13 11.551961
Rsn11_13 sn11_13 sn12_13 11.551961
Rsp11_14 sp11_14 sp12_14 11.551961
Rsn11_14 sn11_14 sn12_14 11.551961
Rsp11_15 sp11_15 sp12_15 11.551961
Rsn11_15 sn11_15 sn12_15 11.551961
Rsp11_16 sp11_16 sp12_16 11.551961
Rsn11_16 sn11_16 sn12_16 11.551961
Rsp11_17 sp11_17 sp12_17 11.551961
Rsn11_17 sn11_17 sn12_17 11.551961
Rsp11_18 sp11_18 sp12_18 11.551961
Rsn11_18 sn11_18 sn12_18 11.551961
Rsp11_19 sp11_19 sp12_19 11.551961
Rsn11_19 sn11_19 sn12_19 11.551961
Rsp11_20 sp11_20 sp12_20 11.551961
Rsn11_20 sn11_20 sn12_20 11.551961
Rsp11_21 sp11_21 sp12_21 11.551961
Rsn11_21 sn11_21 sn12_21 11.551961
Rsp11_22 sp11_22 sp12_22 11.551961
Rsn11_22 sn11_22 sn12_22 11.551961
Rsp11_23 sp11_23 sp12_23 11.551961
Rsn11_23 sn11_23 sn12_23 11.551961
Rsp11_24 sp11_24 sp12_24 11.551961
Rsn11_24 sn11_24 sn12_24 11.551961
Rsp11_25 sp11_25 sp12_25 11.551961
Rsn11_25 sn11_25 sn12_25 11.551961
Rsp11_26 sp11_26 sp12_26 11.551961
Rsn11_26 sn11_26 sn12_26 11.551961
Rsp11_27 sp11_27 sp12_27 11.551961
Rsn11_27 sn11_27 sn12_27 11.551961
Rsp11_28 sp11_28 sp12_28 11.551961
Rsn11_28 sn11_28 sn12_28 11.551961
Rsp11_29 sp11_29 sp12_29 11.551961
Rsn11_29 sn11_29 sn12_29 11.551961
Rsp11_30 sp11_30 sp12_30 11.551961
Rsn11_30 sn11_30 sn12_30 11.551961
Rsp11_31 sp11_31 sp12_31 11.551961
Rsn11_31 sn11_31 sn12_31 11.551961
Rsp11_32 sp11_32 sp12_32 11.551961
Rsn11_32 sn11_32 sn12_32 11.551961
Rsp11_33 sp11_33 sp12_33 11.551961
Rsn11_33 sn11_33 sn12_33 11.551961
Rsp11_34 sp11_34 sp12_34 11.551961
Rsn11_34 sn11_34 sn12_34 11.551961
Rsp11_35 sp11_35 sp12_35 11.551961
Rsn11_35 sn11_35 sn12_35 11.551961
Rsp11_36 sp11_36 sp12_36 11.551961
Rsn11_36 sn11_36 sn12_36 11.551961
Rsp11_37 sp11_37 sp12_37 11.551961
Rsn11_37 sn11_37 sn12_37 11.551961
Rsp11_38 sp11_38 sp12_38 11.551961
Rsn11_38 sn11_38 sn12_38 11.551961
Rsp11_39 sp11_39 sp12_39 11.551961
Rsn11_39 sn11_39 sn12_39 11.551961
Rsp11_40 sp11_40 sp12_40 11.551961
Rsn11_40 sn11_40 sn12_40 11.551961
Rsp11_41 sp11_41 sp12_41 11.551961
Rsn11_41 sn11_41 sn12_41 11.551961
Rsp11_42 sp11_42 sp12_42 11.551961
Rsn11_42 sn11_42 sn12_42 11.551961
Rsp11_43 sp11_43 sp12_43 11.551961
Rsn11_43 sn11_43 sn12_43 11.551961
Rsp11_44 sp11_44 sp12_44 11.551961
Rsn11_44 sn11_44 sn12_44 11.551961
Rsp11_45 sp11_45 sp12_45 11.551961
Rsn11_45 sn11_45 sn12_45 11.551961
Rsp11_46 sp11_46 sp12_46 11.551961
Rsn11_46 sn11_46 sn12_46 11.551961
Rsp11_47 sp11_47 sp12_47 11.551961
Rsn11_47 sn11_47 sn12_47 11.551961
Rsp11_48 sp11_48 sp12_48 11.551961
Rsn11_48 sn11_48 sn12_48 11.551961
Rsp11_49 sp11_49 sp12_49 11.551961
Rsn11_49 sn11_49 sn12_49 11.551961
Rsp11_50 sp11_50 sp12_50 11.551961
Rsn11_50 sn11_50 sn12_50 11.551961
Rsp11_51 sp11_51 sp12_51 11.551961
Rsn11_51 sn11_51 sn12_51 11.551961
Rsp11_52 sp11_52 sp12_52 11.551961
Rsn11_52 sn11_52 sn12_52 11.551961
Rsp11_53 sp11_53 sp12_53 11.551961
Rsn11_53 sn11_53 sn12_53 11.551961
Rsp11_54 sp11_54 sp12_54 11.551961
Rsn11_54 sn11_54 sn12_54 11.551961
Rsp11_55 sp11_55 sp12_55 11.551961
Rsn11_55 sn11_55 sn12_55 11.551961
Rsp11_56 sp11_56 sp12_56 11.551961
Rsn11_56 sn11_56 sn12_56 11.551961
Rsp11_57 sp11_57 sp12_57 11.551961
Rsn11_57 sn11_57 sn12_57 11.551961
Rsp11_58 sp11_58 sp12_58 11.551961
Rsn11_58 sn11_58 sn12_58 11.551961
Rsp11_59 sp11_59 sp12_59 11.551961
Rsn11_59 sn11_59 sn12_59 11.551961
Rsp11_60 sp11_60 sp12_60 11.551961
Rsn11_60 sn11_60 sn12_60 11.551961
Rsp11_61 sp11_61 sp12_61 11.551961
Rsn11_61 sn11_61 sn12_61 11.551961
Rsp11_62 sp11_62 sp12_62 11.551961
Rsn11_62 sn11_62 sn12_62 11.551961
Rsp11_63 sp11_63 sp12_63 11.551961
Rsn11_63 sn11_63 sn12_63 11.551961
Rsp11_64 sp11_64 sp12_64 11.551961
Rsn11_64 sn11_64 sn12_64 11.551961
Rsp11_65 sp11_65 sp12_65 11.551961
Rsn11_65 sn11_65 sn12_65 11.551961
Rsp11_66 sp11_66 sp12_66 11.551961
Rsn11_66 sn11_66 sn12_66 11.551961
Rsp11_67 sp11_67 sp12_67 11.551961
Rsn11_67 sn11_67 sn12_67 11.551961
Rsp11_68 sp11_68 sp12_68 11.551961
Rsn11_68 sn11_68 sn12_68 11.551961
Rsp11_69 sp11_69 sp12_69 11.551961
Rsn11_69 sn11_69 sn12_69 11.551961
Rsp11_70 sp11_70 sp12_70 11.551961
Rsn11_70 sn11_70 sn12_70 11.551961
Rsp11_71 sp11_71 sp12_71 11.551961
Rsn11_71 sn11_71 sn12_71 11.551961
Rsp11_72 sp11_72 sp12_72 11.551961
Rsn11_72 sn11_72 sn12_72 11.551961
Rsp11_73 sp11_73 sp12_73 11.551961
Rsn11_73 sn11_73 sn12_73 11.551961
Rsp11_74 sp11_74 sp12_74 11.551961
Rsn11_74 sn11_74 sn12_74 11.551961
Rsp11_75 sp11_75 sp12_75 11.551961
Rsn11_75 sn11_75 sn12_75 11.551961
Rsp11_76 sp11_76 sp12_76 11.551961
Rsn11_76 sn11_76 sn12_76 11.551961
Rsp11_77 sp11_77 sp12_77 11.551961
Rsn11_77 sn11_77 sn12_77 11.551961
Rsp11_78 sp11_78 sp12_78 11.551961
Rsn11_78 sn11_78 sn12_78 11.551961
Rsp11_79 sp11_79 sp12_79 11.551961
Rsn11_79 sn11_79 sn12_79 11.551961
Rsp11_80 sp11_80 sp12_80 11.551961
Rsn11_80 sn11_80 sn12_80 11.551961
Rsp11_81 sp11_81 sp12_81 11.551961
Rsn11_81 sn11_81 sn12_81 11.551961
Rsp11_82 sp11_82 sp12_82 11.551961
Rsn11_82 sn11_82 sn12_82 11.551961
Rsp11_83 sp11_83 sp12_83 11.551961
Rsn11_83 sn11_83 sn12_83 11.551961
Rsp11_84 sp11_84 sp12_84 11.551961
Rsn11_84 sn11_84 sn12_84 11.551961
Rsp12_1 sp12_1 sp13_1 11.551961
Rsn12_1 sn12_1 sn13_1 11.551961
Rsp12_2 sp12_2 sp13_2 11.551961
Rsn12_2 sn12_2 sn13_2 11.551961
Rsp12_3 sp12_3 sp13_3 11.551961
Rsn12_3 sn12_3 sn13_3 11.551961
Rsp12_4 sp12_4 sp13_4 11.551961
Rsn12_4 sn12_4 sn13_4 11.551961
Rsp12_5 sp12_5 sp13_5 11.551961
Rsn12_5 sn12_5 sn13_5 11.551961
Rsp12_6 sp12_6 sp13_6 11.551961
Rsn12_6 sn12_6 sn13_6 11.551961
Rsp12_7 sp12_7 sp13_7 11.551961
Rsn12_7 sn12_7 sn13_7 11.551961
Rsp12_8 sp12_8 sp13_8 11.551961
Rsn12_8 sn12_8 sn13_8 11.551961
Rsp12_9 sp12_9 sp13_9 11.551961
Rsn12_9 sn12_9 sn13_9 11.551961
Rsp12_10 sp12_10 sp13_10 11.551961
Rsn12_10 sn12_10 sn13_10 11.551961
Rsp12_11 sp12_11 sp13_11 11.551961
Rsn12_11 sn12_11 sn13_11 11.551961
Rsp12_12 sp12_12 sp13_12 11.551961
Rsn12_12 sn12_12 sn13_12 11.551961
Rsp12_13 sp12_13 sp13_13 11.551961
Rsn12_13 sn12_13 sn13_13 11.551961
Rsp12_14 sp12_14 sp13_14 11.551961
Rsn12_14 sn12_14 sn13_14 11.551961
Rsp12_15 sp12_15 sp13_15 11.551961
Rsn12_15 sn12_15 sn13_15 11.551961
Rsp12_16 sp12_16 sp13_16 11.551961
Rsn12_16 sn12_16 sn13_16 11.551961
Rsp12_17 sp12_17 sp13_17 11.551961
Rsn12_17 sn12_17 sn13_17 11.551961
Rsp12_18 sp12_18 sp13_18 11.551961
Rsn12_18 sn12_18 sn13_18 11.551961
Rsp12_19 sp12_19 sp13_19 11.551961
Rsn12_19 sn12_19 sn13_19 11.551961
Rsp12_20 sp12_20 sp13_20 11.551961
Rsn12_20 sn12_20 sn13_20 11.551961
Rsp12_21 sp12_21 sp13_21 11.551961
Rsn12_21 sn12_21 sn13_21 11.551961
Rsp12_22 sp12_22 sp13_22 11.551961
Rsn12_22 sn12_22 sn13_22 11.551961
Rsp12_23 sp12_23 sp13_23 11.551961
Rsn12_23 sn12_23 sn13_23 11.551961
Rsp12_24 sp12_24 sp13_24 11.551961
Rsn12_24 sn12_24 sn13_24 11.551961
Rsp12_25 sp12_25 sp13_25 11.551961
Rsn12_25 sn12_25 sn13_25 11.551961
Rsp12_26 sp12_26 sp13_26 11.551961
Rsn12_26 sn12_26 sn13_26 11.551961
Rsp12_27 sp12_27 sp13_27 11.551961
Rsn12_27 sn12_27 sn13_27 11.551961
Rsp12_28 sp12_28 sp13_28 11.551961
Rsn12_28 sn12_28 sn13_28 11.551961
Rsp12_29 sp12_29 sp13_29 11.551961
Rsn12_29 sn12_29 sn13_29 11.551961
Rsp12_30 sp12_30 sp13_30 11.551961
Rsn12_30 sn12_30 sn13_30 11.551961
Rsp12_31 sp12_31 sp13_31 11.551961
Rsn12_31 sn12_31 sn13_31 11.551961
Rsp12_32 sp12_32 sp13_32 11.551961
Rsn12_32 sn12_32 sn13_32 11.551961
Rsp12_33 sp12_33 sp13_33 11.551961
Rsn12_33 sn12_33 sn13_33 11.551961
Rsp12_34 sp12_34 sp13_34 11.551961
Rsn12_34 sn12_34 sn13_34 11.551961
Rsp12_35 sp12_35 sp13_35 11.551961
Rsn12_35 sn12_35 sn13_35 11.551961
Rsp12_36 sp12_36 sp13_36 11.551961
Rsn12_36 sn12_36 sn13_36 11.551961
Rsp12_37 sp12_37 sp13_37 11.551961
Rsn12_37 sn12_37 sn13_37 11.551961
Rsp12_38 sp12_38 sp13_38 11.551961
Rsn12_38 sn12_38 sn13_38 11.551961
Rsp12_39 sp12_39 sp13_39 11.551961
Rsn12_39 sn12_39 sn13_39 11.551961
Rsp12_40 sp12_40 sp13_40 11.551961
Rsn12_40 sn12_40 sn13_40 11.551961
Rsp12_41 sp12_41 sp13_41 11.551961
Rsn12_41 sn12_41 sn13_41 11.551961
Rsp12_42 sp12_42 sp13_42 11.551961
Rsn12_42 sn12_42 sn13_42 11.551961
Rsp12_43 sp12_43 sp13_43 11.551961
Rsn12_43 sn12_43 sn13_43 11.551961
Rsp12_44 sp12_44 sp13_44 11.551961
Rsn12_44 sn12_44 sn13_44 11.551961
Rsp12_45 sp12_45 sp13_45 11.551961
Rsn12_45 sn12_45 sn13_45 11.551961
Rsp12_46 sp12_46 sp13_46 11.551961
Rsn12_46 sn12_46 sn13_46 11.551961
Rsp12_47 sp12_47 sp13_47 11.551961
Rsn12_47 sn12_47 sn13_47 11.551961
Rsp12_48 sp12_48 sp13_48 11.551961
Rsn12_48 sn12_48 sn13_48 11.551961
Rsp12_49 sp12_49 sp13_49 11.551961
Rsn12_49 sn12_49 sn13_49 11.551961
Rsp12_50 sp12_50 sp13_50 11.551961
Rsn12_50 sn12_50 sn13_50 11.551961
Rsp12_51 sp12_51 sp13_51 11.551961
Rsn12_51 sn12_51 sn13_51 11.551961
Rsp12_52 sp12_52 sp13_52 11.551961
Rsn12_52 sn12_52 sn13_52 11.551961
Rsp12_53 sp12_53 sp13_53 11.551961
Rsn12_53 sn12_53 sn13_53 11.551961
Rsp12_54 sp12_54 sp13_54 11.551961
Rsn12_54 sn12_54 sn13_54 11.551961
Rsp12_55 sp12_55 sp13_55 11.551961
Rsn12_55 sn12_55 sn13_55 11.551961
Rsp12_56 sp12_56 sp13_56 11.551961
Rsn12_56 sn12_56 sn13_56 11.551961
Rsp12_57 sp12_57 sp13_57 11.551961
Rsn12_57 sn12_57 sn13_57 11.551961
Rsp12_58 sp12_58 sp13_58 11.551961
Rsn12_58 sn12_58 sn13_58 11.551961
Rsp12_59 sp12_59 sp13_59 11.551961
Rsn12_59 sn12_59 sn13_59 11.551961
Rsp12_60 sp12_60 sp13_60 11.551961
Rsn12_60 sn12_60 sn13_60 11.551961
Rsp12_61 sp12_61 sp13_61 11.551961
Rsn12_61 sn12_61 sn13_61 11.551961
Rsp12_62 sp12_62 sp13_62 11.551961
Rsn12_62 sn12_62 sn13_62 11.551961
Rsp12_63 sp12_63 sp13_63 11.551961
Rsn12_63 sn12_63 sn13_63 11.551961
Rsp12_64 sp12_64 sp13_64 11.551961
Rsn12_64 sn12_64 sn13_64 11.551961
Rsp12_65 sp12_65 sp13_65 11.551961
Rsn12_65 sn12_65 sn13_65 11.551961
Rsp12_66 sp12_66 sp13_66 11.551961
Rsn12_66 sn12_66 sn13_66 11.551961
Rsp12_67 sp12_67 sp13_67 11.551961
Rsn12_67 sn12_67 sn13_67 11.551961
Rsp12_68 sp12_68 sp13_68 11.551961
Rsn12_68 sn12_68 sn13_68 11.551961
Rsp12_69 sp12_69 sp13_69 11.551961
Rsn12_69 sn12_69 sn13_69 11.551961
Rsp12_70 sp12_70 sp13_70 11.551961
Rsn12_70 sn12_70 sn13_70 11.551961
Rsp12_71 sp12_71 sp13_71 11.551961
Rsn12_71 sn12_71 sn13_71 11.551961
Rsp12_72 sp12_72 sp13_72 11.551961
Rsn12_72 sn12_72 sn13_72 11.551961
Rsp12_73 sp12_73 sp13_73 11.551961
Rsn12_73 sn12_73 sn13_73 11.551961
Rsp12_74 sp12_74 sp13_74 11.551961
Rsn12_74 sn12_74 sn13_74 11.551961
Rsp12_75 sp12_75 sp13_75 11.551961
Rsn12_75 sn12_75 sn13_75 11.551961
Rsp12_76 sp12_76 sp13_76 11.551961
Rsn12_76 sn12_76 sn13_76 11.551961
Rsp12_77 sp12_77 sp13_77 11.551961
Rsn12_77 sn12_77 sn13_77 11.551961
Rsp12_78 sp12_78 sp13_78 11.551961
Rsn12_78 sn12_78 sn13_78 11.551961
Rsp12_79 sp12_79 sp13_79 11.551961
Rsn12_79 sn12_79 sn13_79 11.551961
Rsp12_80 sp12_80 sp13_80 11.551961
Rsn12_80 sn12_80 sn13_80 11.551961
Rsp12_81 sp12_81 sp13_81 11.551961
Rsn12_81 sn12_81 sn13_81 11.551961
Rsp12_82 sp12_82 sp13_82 11.551961
Rsn12_82 sn12_82 sn13_82 11.551961
Rsp12_83 sp12_83 sp13_83 11.551961
Rsn12_83 sn12_83 sn13_83 11.551961
Rsp12_84 sp12_84 sp13_84 11.551961
Rsn12_84 sn12_84 sn13_84 11.551961
Rsp13_1 sp13_1 sp14_1 11.551961
Rsn13_1 sn13_1 sn14_1 11.551961
Rsp13_2 sp13_2 sp14_2 11.551961
Rsn13_2 sn13_2 sn14_2 11.551961
Rsp13_3 sp13_3 sp14_3 11.551961
Rsn13_3 sn13_3 sn14_3 11.551961
Rsp13_4 sp13_4 sp14_4 11.551961
Rsn13_4 sn13_4 sn14_4 11.551961
Rsp13_5 sp13_5 sp14_5 11.551961
Rsn13_5 sn13_5 sn14_5 11.551961
Rsp13_6 sp13_6 sp14_6 11.551961
Rsn13_6 sn13_6 sn14_6 11.551961
Rsp13_7 sp13_7 sp14_7 11.551961
Rsn13_7 sn13_7 sn14_7 11.551961
Rsp13_8 sp13_8 sp14_8 11.551961
Rsn13_8 sn13_8 sn14_8 11.551961
Rsp13_9 sp13_9 sp14_9 11.551961
Rsn13_9 sn13_9 sn14_9 11.551961
Rsp13_10 sp13_10 sp14_10 11.551961
Rsn13_10 sn13_10 sn14_10 11.551961
Rsp13_11 sp13_11 sp14_11 11.551961
Rsn13_11 sn13_11 sn14_11 11.551961
Rsp13_12 sp13_12 sp14_12 11.551961
Rsn13_12 sn13_12 sn14_12 11.551961
Rsp13_13 sp13_13 sp14_13 11.551961
Rsn13_13 sn13_13 sn14_13 11.551961
Rsp13_14 sp13_14 sp14_14 11.551961
Rsn13_14 sn13_14 sn14_14 11.551961
Rsp13_15 sp13_15 sp14_15 11.551961
Rsn13_15 sn13_15 sn14_15 11.551961
Rsp13_16 sp13_16 sp14_16 11.551961
Rsn13_16 sn13_16 sn14_16 11.551961
Rsp13_17 sp13_17 sp14_17 11.551961
Rsn13_17 sn13_17 sn14_17 11.551961
Rsp13_18 sp13_18 sp14_18 11.551961
Rsn13_18 sn13_18 sn14_18 11.551961
Rsp13_19 sp13_19 sp14_19 11.551961
Rsn13_19 sn13_19 sn14_19 11.551961
Rsp13_20 sp13_20 sp14_20 11.551961
Rsn13_20 sn13_20 sn14_20 11.551961
Rsp13_21 sp13_21 sp14_21 11.551961
Rsn13_21 sn13_21 sn14_21 11.551961
Rsp13_22 sp13_22 sp14_22 11.551961
Rsn13_22 sn13_22 sn14_22 11.551961
Rsp13_23 sp13_23 sp14_23 11.551961
Rsn13_23 sn13_23 sn14_23 11.551961
Rsp13_24 sp13_24 sp14_24 11.551961
Rsn13_24 sn13_24 sn14_24 11.551961
Rsp13_25 sp13_25 sp14_25 11.551961
Rsn13_25 sn13_25 sn14_25 11.551961
Rsp13_26 sp13_26 sp14_26 11.551961
Rsn13_26 sn13_26 sn14_26 11.551961
Rsp13_27 sp13_27 sp14_27 11.551961
Rsn13_27 sn13_27 sn14_27 11.551961
Rsp13_28 sp13_28 sp14_28 11.551961
Rsn13_28 sn13_28 sn14_28 11.551961
Rsp13_29 sp13_29 sp14_29 11.551961
Rsn13_29 sn13_29 sn14_29 11.551961
Rsp13_30 sp13_30 sp14_30 11.551961
Rsn13_30 sn13_30 sn14_30 11.551961
Rsp13_31 sp13_31 sp14_31 11.551961
Rsn13_31 sn13_31 sn14_31 11.551961
Rsp13_32 sp13_32 sp14_32 11.551961
Rsn13_32 sn13_32 sn14_32 11.551961
Rsp13_33 sp13_33 sp14_33 11.551961
Rsn13_33 sn13_33 sn14_33 11.551961
Rsp13_34 sp13_34 sp14_34 11.551961
Rsn13_34 sn13_34 sn14_34 11.551961
Rsp13_35 sp13_35 sp14_35 11.551961
Rsn13_35 sn13_35 sn14_35 11.551961
Rsp13_36 sp13_36 sp14_36 11.551961
Rsn13_36 sn13_36 sn14_36 11.551961
Rsp13_37 sp13_37 sp14_37 11.551961
Rsn13_37 sn13_37 sn14_37 11.551961
Rsp13_38 sp13_38 sp14_38 11.551961
Rsn13_38 sn13_38 sn14_38 11.551961
Rsp13_39 sp13_39 sp14_39 11.551961
Rsn13_39 sn13_39 sn14_39 11.551961
Rsp13_40 sp13_40 sp14_40 11.551961
Rsn13_40 sn13_40 sn14_40 11.551961
Rsp13_41 sp13_41 sp14_41 11.551961
Rsn13_41 sn13_41 sn14_41 11.551961
Rsp13_42 sp13_42 sp14_42 11.551961
Rsn13_42 sn13_42 sn14_42 11.551961
Rsp13_43 sp13_43 sp14_43 11.551961
Rsn13_43 sn13_43 sn14_43 11.551961
Rsp13_44 sp13_44 sp14_44 11.551961
Rsn13_44 sn13_44 sn14_44 11.551961
Rsp13_45 sp13_45 sp14_45 11.551961
Rsn13_45 sn13_45 sn14_45 11.551961
Rsp13_46 sp13_46 sp14_46 11.551961
Rsn13_46 sn13_46 sn14_46 11.551961
Rsp13_47 sp13_47 sp14_47 11.551961
Rsn13_47 sn13_47 sn14_47 11.551961
Rsp13_48 sp13_48 sp14_48 11.551961
Rsn13_48 sn13_48 sn14_48 11.551961
Rsp13_49 sp13_49 sp14_49 11.551961
Rsn13_49 sn13_49 sn14_49 11.551961
Rsp13_50 sp13_50 sp14_50 11.551961
Rsn13_50 sn13_50 sn14_50 11.551961
Rsp13_51 sp13_51 sp14_51 11.551961
Rsn13_51 sn13_51 sn14_51 11.551961
Rsp13_52 sp13_52 sp14_52 11.551961
Rsn13_52 sn13_52 sn14_52 11.551961
Rsp13_53 sp13_53 sp14_53 11.551961
Rsn13_53 sn13_53 sn14_53 11.551961
Rsp13_54 sp13_54 sp14_54 11.551961
Rsn13_54 sn13_54 sn14_54 11.551961
Rsp13_55 sp13_55 sp14_55 11.551961
Rsn13_55 sn13_55 sn14_55 11.551961
Rsp13_56 sp13_56 sp14_56 11.551961
Rsn13_56 sn13_56 sn14_56 11.551961
Rsp13_57 sp13_57 sp14_57 11.551961
Rsn13_57 sn13_57 sn14_57 11.551961
Rsp13_58 sp13_58 sp14_58 11.551961
Rsn13_58 sn13_58 sn14_58 11.551961
Rsp13_59 sp13_59 sp14_59 11.551961
Rsn13_59 sn13_59 sn14_59 11.551961
Rsp13_60 sp13_60 sp14_60 11.551961
Rsn13_60 sn13_60 sn14_60 11.551961
Rsp13_61 sp13_61 sp14_61 11.551961
Rsn13_61 sn13_61 sn14_61 11.551961
Rsp13_62 sp13_62 sp14_62 11.551961
Rsn13_62 sn13_62 sn14_62 11.551961
Rsp13_63 sp13_63 sp14_63 11.551961
Rsn13_63 sn13_63 sn14_63 11.551961
Rsp13_64 sp13_64 sp14_64 11.551961
Rsn13_64 sn13_64 sn14_64 11.551961
Rsp13_65 sp13_65 sp14_65 11.551961
Rsn13_65 sn13_65 sn14_65 11.551961
Rsp13_66 sp13_66 sp14_66 11.551961
Rsn13_66 sn13_66 sn14_66 11.551961
Rsp13_67 sp13_67 sp14_67 11.551961
Rsn13_67 sn13_67 sn14_67 11.551961
Rsp13_68 sp13_68 sp14_68 11.551961
Rsn13_68 sn13_68 sn14_68 11.551961
Rsp13_69 sp13_69 sp14_69 11.551961
Rsn13_69 sn13_69 sn14_69 11.551961
Rsp13_70 sp13_70 sp14_70 11.551961
Rsn13_70 sn13_70 sn14_70 11.551961
Rsp13_71 sp13_71 sp14_71 11.551961
Rsn13_71 sn13_71 sn14_71 11.551961
Rsp13_72 sp13_72 sp14_72 11.551961
Rsn13_72 sn13_72 sn14_72 11.551961
Rsp13_73 sp13_73 sp14_73 11.551961
Rsn13_73 sn13_73 sn14_73 11.551961
Rsp13_74 sp13_74 sp14_74 11.551961
Rsn13_74 sn13_74 sn14_74 11.551961
Rsp13_75 sp13_75 sp14_75 11.551961
Rsn13_75 sn13_75 sn14_75 11.551961
Rsp13_76 sp13_76 sp14_76 11.551961
Rsn13_76 sn13_76 sn14_76 11.551961
Rsp13_77 sp13_77 sp14_77 11.551961
Rsn13_77 sn13_77 sn14_77 11.551961
Rsp13_78 sp13_78 sp14_78 11.551961
Rsn13_78 sn13_78 sn14_78 11.551961
Rsp13_79 sp13_79 sp14_79 11.551961
Rsn13_79 sn13_79 sn14_79 11.551961
Rsp13_80 sp13_80 sp14_80 11.551961
Rsn13_80 sn13_80 sn14_80 11.551961
Rsp13_81 sp13_81 sp14_81 11.551961
Rsn13_81 sn13_81 sn14_81 11.551961
Rsp13_82 sp13_82 sp14_82 11.551961
Rsn13_82 sn13_82 sn14_82 11.551961
Rsp13_83 sp13_83 sp14_83 11.551961
Rsn13_83 sn13_83 sn14_83 11.551961
Rsp13_84 sp13_84 sp14_84 11.551961
Rsn13_84 sn13_84 sn14_84 11.551961
Rsp14_1 sp14_1 sp15_1 11.551961
Rsn14_1 sn14_1 sn15_1 11.551961
Rsp14_2 sp14_2 sp15_2 11.551961
Rsn14_2 sn14_2 sn15_2 11.551961
Rsp14_3 sp14_3 sp15_3 11.551961
Rsn14_3 sn14_3 sn15_3 11.551961
Rsp14_4 sp14_4 sp15_4 11.551961
Rsn14_4 sn14_4 sn15_4 11.551961
Rsp14_5 sp14_5 sp15_5 11.551961
Rsn14_5 sn14_5 sn15_5 11.551961
Rsp14_6 sp14_6 sp15_6 11.551961
Rsn14_6 sn14_6 sn15_6 11.551961
Rsp14_7 sp14_7 sp15_7 11.551961
Rsn14_7 sn14_7 sn15_7 11.551961
Rsp14_8 sp14_8 sp15_8 11.551961
Rsn14_8 sn14_8 sn15_8 11.551961
Rsp14_9 sp14_9 sp15_9 11.551961
Rsn14_9 sn14_9 sn15_9 11.551961
Rsp14_10 sp14_10 sp15_10 11.551961
Rsn14_10 sn14_10 sn15_10 11.551961
Rsp14_11 sp14_11 sp15_11 11.551961
Rsn14_11 sn14_11 sn15_11 11.551961
Rsp14_12 sp14_12 sp15_12 11.551961
Rsn14_12 sn14_12 sn15_12 11.551961
Rsp14_13 sp14_13 sp15_13 11.551961
Rsn14_13 sn14_13 sn15_13 11.551961
Rsp14_14 sp14_14 sp15_14 11.551961
Rsn14_14 sn14_14 sn15_14 11.551961
Rsp14_15 sp14_15 sp15_15 11.551961
Rsn14_15 sn14_15 sn15_15 11.551961
Rsp14_16 sp14_16 sp15_16 11.551961
Rsn14_16 sn14_16 sn15_16 11.551961
Rsp14_17 sp14_17 sp15_17 11.551961
Rsn14_17 sn14_17 sn15_17 11.551961
Rsp14_18 sp14_18 sp15_18 11.551961
Rsn14_18 sn14_18 sn15_18 11.551961
Rsp14_19 sp14_19 sp15_19 11.551961
Rsn14_19 sn14_19 sn15_19 11.551961
Rsp14_20 sp14_20 sp15_20 11.551961
Rsn14_20 sn14_20 sn15_20 11.551961
Rsp14_21 sp14_21 sp15_21 11.551961
Rsn14_21 sn14_21 sn15_21 11.551961
Rsp14_22 sp14_22 sp15_22 11.551961
Rsn14_22 sn14_22 sn15_22 11.551961
Rsp14_23 sp14_23 sp15_23 11.551961
Rsn14_23 sn14_23 sn15_23 11.551961
Rsp14_24 sp14_24 sp15_24 11.551961
Rsn14_24 sn14_24 sn15_24 11.551961
Rsp14_25 sp14_25 sp15_25 11.551961
Rsn14_25 sn14_25 sn15_25 11.551961
Rsp14_26 sp14_26 sp15_26 11.551961
Rsn14_26 sn14_26 sn15_26 11.551961
Rsp14_27 sp14_27 sp15_27 11.551961
Rsn14_27 sn14_27 sn15_27 11.551961
Rsp14_28 sp14_28 sp15_28 11.551961
Rsn14_28 sn14_28 sn15_28 11.551961
Rsp14_29 sp14_29 sp15_29 11.551961
Rsn14_29 sn14_29 sn15_29 11.551961
Rsp14_30 sp14_30 sp15_30 11.551961
Rsn14_30 sn14_30 sn15_30 11.551961
Rsp14_31 sp14_31 sp15_31 11.551961
Rsn14_31 sn14_31 sn15_31 11.551961
Rsp14_32 sp14_32 sp15_32 11.551961
Rsn14_32 sn14_32 sn15_32 11.551961
Rsp14_33 sp14_33 sp15_33 11.551961
Rsn14_33 sn14_33 sn15_33 11.551961
Rsp14_34 sp14_34 sp15_34 11.551961
Rsn14_34 sn14_34 sn15_34 11.551961
Rsp14_35 sp14_35 sp15_35 11.551961
Rsn14_35 sn14_35 sn15_35 11.551961
Rsp14_36 sp14_36 sp15_36 11.551961
Rsn14_36 sn14_36 sn15_36 11.551961
Rsp14_37 sp14_37 sp15_37 11.551961
Rsn14_37 sn14_37 sn15_37 11.551961
Rsp14_38 sp14_38 sp15_38 11.551961
Rsn14_38 sn14_38 sn15_38 11.551961
Rsp14_39 sp14_39 sp15_39 11.551961
Rsn14_39 sn14_39 sn15_39 11.551961
Rsp14_40 sp14_40 sp15_40 11.551961
Rsn14_40 sn14_40 sn15_40 11.551961
Rsp14_41 sp14_41 sp15_41 11.551961
Rsn14_41 sn14_41 sn15_41 11.551961
Rsp14_42 sp14_42 sp15_42 11.551961
Rsn14_42 sn14_42 sn15_42 11.551961
Rsp14_43 sp14_43 sp15_43 11.551961
Rsn14_43 sn14_43 sn15_43 11.551961
Rsp14_44 sp14_44 sp15_44 11.551961
Rsn14_44 sn14_44 sn15_44 11.551961
Rsp14_45 sp14_45 sp15_45 11.551961
Rsn14_45 sn14_45 sn15_45 11.551961
Rsp14_46 sp14_46 sp15_46 11.551961
Rsn14_46 sn14_46 sn15_46 11.551961
Rsp14_47 sp14_47 sp15_47 11.551961
Rsn14_47 sn14_47 sn15_47 11.551961
Rsp14_48 sp14_48 sp15_48 11.551961
Rsn14_48 sn14_48 sn15_48 11.551961
Rsp14_49 sp14_49 sp15_49 11.551961
Rsn14_49 sn14_49 sn15_49 11.551961
Rsp14_50 sp14_50 sp15_50 11.551961
Rsn14_50 sn14_50 sn15_50 11.551961
Rsp14_51 sp14_51 sp15_51 11.551961
Rsn14_51 sn14_51 sn15_51 11.551961
Rsp14_52 sp14_52 sp15_52 11.551961
Rsn14_52 sn14_52 sn15_52 11.551961
Rsp14_53 sp14_53 sp15_53 11.551961
Rsn14_53 sn14_53 sn15_53 11.551961
Rsp14_54 sp14_54 sp15_54 11.551961
Rsn14_54 sn14_54 sn15_54 11.551961
Rsp14_55 sp14_55 sp15_55 11.551961
Rsn14_55 sn14_55 sn15_55 11.551961
Rsp14_56 sp14_56 sp15_56 11.551961
Rsn14_56 sn14_56 sn15_56 11.551961
Rsp14_57 sp14_57 sp15_57 11.551961
Rsn14_57 sn14_57 sn15_57 11.551961
Rsp14_58 sp14_58 sp15_58 11.551961
Rsn14_58 sn14_58 sn15_58 11.551961
Rsp14_59 sp14_59 sp15_59 11.551961
Rsn14_59 sn14_59 sn15_59 11.551961
Rsp14_60 sp14_60 sp15_60 11.551961
Rsn14_60 sn14_60 sn15_60 11.551961
Rsp14_61 sp14_61 sp15_61 11.551961
Rsn14_61 sn14_61 sn15_61 11.551961
Rsp14_62 sp14_62 sp15_62 11.551961
Rsn14_62 sn14_62 sn15_62 11.551961
Rsp14_63 sp14_63 sp15_63 11.551961
Rsn14_63 sn14_63 sn15_63 11.551961
Rsp14_64 sp14_64 sp15_64 11.551961
Rsn14_64 sn14_64 sn15_64 11.551961
Rsp14_65 sp14_65 sp15_65 11.551961
Rsn14_65 sn14_65 sn15_65 11.551961
Rsp14_66 sp14_66 sp15_66 11.551961
Rsn14_66 sn14_66 sn15_66 11.551961
Rsp14_67 sp14_67 sp15_67 11.551961
Rsn14_67 sn14_67 sn15_67 11.551961
Rsp14_68 sp14_68 sp15_68 11.551961
Rsn14_68 sn14_68 sn15_68 11.551961
Rsp14_69 sp14_69 sp15_69 11.551961
Rsn14_69 sn14_69 sn15_69 11.551961
Rsp14_70 sp14_70 sp15_70 11.551961
Rsn14_70 sn14_70 sn15_70 11.551961
Rsp14_71 sp14_71 sp15_71 11.551961
Rsn14_71 sn14_71 sn15_71 11.551961
Rsp14_72 sp14_72 sp15_72 11.551961
Rsn14_72 sn14_72 sn15_72 11.551961
Rsp14_73 sp14_73 sp15_73 11.551961
Rsn14_73 sn14_73 sn15_73 11.551961
Rsp14_74 sp14_74 sp15_74 11.551961
Rsn14_74 sn14_74 sn15_74 11.551961
Rsp14_75 sp14_75 sp15_75 11.551961
Rsn14_75 sn14_75 sn15_75 11.551961
Rsp14_76 sp14_76 sp15_76 11.551961
Rsn14_76 sn14_76 sn15_76 11.551961
Rsp14_77 sp14_77 sp15_77 11.551961
Rsn14_77 sn14_77 sn15_77 11.551961
Rsp14_78 sp14_78 sp15_78 11.551961
Rsn14_78 sn14_78 sn15_78 11.551961
Rsp14_79 sp14_79 sp15_79 11.551961
Rsn14_79 sn14_79 sn15_79 11.551961
Rsp14_80 sp14_80 sp15_80 11.551961
Rsn14_80 sn14_80 sn15_80 11.551961
Rsp14_81 sp14_81 sp15_81 11.551961
Rsn14_81 sn14_81 sn15_81 11.551961
Rsp14_82 sp14_82 sp15_82 11.551961
Rsn14_82 sn14_82 sn15_82 11.551961
Rsp14_83 sp14_83 sp15_83 11.551961
Rsn14_83 sn14_83 sn15_83 11.551961
Rsp14_84 sp14_84 sp15_84 11.551961
Rsn14_84 sn14_84 sn15_84 11.551961
Rsp15_1 sp15_1 sp16_1 11.551961
Rsn15_1 sn15_1 sn16_1 11.551961
Rsp15_2 sp15_2 sp16_2 11.551961
Rsn15_2 sn15_2 sn16_2 11.551961
Rsp15_3 sp15_3 sp16_3 11.551961
Rsn15_3 sn15_3 sn16_3 11.551961
Rsp15_4 sp15_4 sp16_4 11.551961
Rsn15_4 sn15_4 sn16_4 11.551961
Rsp15_5 sp15_5 sp16_5 11.551961
Rsn15_5 sn15_5 sn16_5 11.551961
Rsp15_6 sp15_6 sp16_6 11.551961
Rsn15_6 sn15_6 sn16_6 11.551961
Rsp15_7 sp15_7 sp16_7 11.551961
Rsn15_7 sn15_7 sn16_7 11.551961
Rsp15_8 sp15_8 sp16_8 11.551961
Rsn15_8 sn15_8 sn16_8 11.551961
Rsp15_9 sp15_9 sp16_9 11.551961
Rsn15_9 sn15_9 sn16_9 11.551961
Rsp15_10 sp15_10 sp16_10 11.551961
Rsn15_10 sn15_10 sn16_10 11.551961
Rsp15_11 sp15_11 sp16_11 11.551961
Rsn15_11 sn15_11 sn16_11 11.551961
Rsp15_12 sp15_12 sp16_12 11.551961
Rsn15_12 sn15_12 sn16_12 11.551961
Rsp15_13 sp15_13 sp16_13 11.551961
Rsn15_13 sn15_13 sn16_13 11.551961
Rsp15_14 sp15_14 sp16_14 11.551961
Rsn15_14 sn15_14 sn16_14 11.551961
Rsp15_15 sp15_15 sp16_15 11.551961
Rsn15_15 sn15_15 sn16_15 11.551961
Rsp15_16 sp15_16 sp16_16 11.551961
Rsn15_16 sn15_16 sn16_16 11.551961
Rsp15_17 sp15_17 sp16_17 11.551961
Rsn15_17 sn15_17 sn16_17 11.551961
Rsp15_18 sp15_18 sp16_18 11.551961
Rsn15_18 sn15_18 sn16_18 11.551961
Rsp15_19 sp15_19 sp16_19 11.551961
Rsn15_19 sn15_19 sn16_19 11.551961
Rsp15_20 sp15_20 sp16_20 11.551961
Rsn15_20 sn15_20 sn16_20 11.551961
Rsp15_21 sp15_21 sp16_21 11.551961
Rsn15_21 sn15_21 sn16_21 11.551961
Rsp15_22 sp15_22 sp16_22 11.551961
Rsn15_22 sn15_22 sn16_22 11.551961
Rsp15_23 sp15_23 sp16_23 11.551961
Rsn15_23 sn15_23 sn16_23 11.551961
Rsp15_24 sp15_24 sp16_24 11.551961
Rsn15_24 sn15_24 sn16_24 11.551961
Rsp15_25 sp15_25 sp16_25 11.551961
Rsn15_25 sn15_25 sn16_25 11.551961
Rsp15_26 sp15_26 sp16_26 11.551961
Rsn15_26 sn15_26 sn16_26 11.551961
Rsp15_27 sp15_27 sp16_27 11.551961
Rsn15_27 sn15_27 sn16_27 11.551961
Rsp15_28 sp15_28 sp16_28 11.551961
Rsn15_28 sn15_28 sn16_28 11.551961
Rsp15_29 sp15_29 sp16_29 11.551961
Rsn15_29 sn15_29 sn16_29 11.551961
Rsp15_30 sp15_30 sp16_30 11.551961
Rsn15_30 sn15_30 sn16_30 11.551961
Rsp15_31 sp15_31 sp16_31 11.551961
Rsn15_31 sn15_31 sn16_31 11.551961
Rsp15_32 sp15_32 sp16_32 11.551961
Rsn15_32 sn15_32 sn16_32 11.551961
Rsp15_33 sp15_33 sp16_33 11.551961
Rsn15_33 sn15_33 sn16_33 11.551961
Rsp15_34 sp15_34 sp16_34 11.551961
Rsn15_34 sn15_34 sn16_34 11.551961
Rsp15_35 sp15_35 sp16_35 11.551961
Rsn15_35 sn15_35 sn16_35 11.551961
Rsp15_36 sp15_36 sp16_36 11.551961
Rsn15_36 sn15_36 sn16_36 11.551961
Rsp15_37 sp15_37 sp16_37 11.551961
Rsn15_37 sn15_37 sn16_37 11.551961
Rsp15_38 sp15_38 sp16_38 11.551961
Rsn15_38 sn15_38 sn16_38 11.551961
Rsp15_39 sp15_39 sp16_39 11.551961
Rsn15_39 sn15_39 sn16_39 11.551961
Rsp15_40 sp15_40 sp16_40 11.551961
Rsn15_40 sn15_40 sn16_40 11.551961
Rsp15_41 sp15_41 sp16_41 11.551961
Rsn15_41 sn15_41 sn16_41 11.551961
Rsp15_42 sp15_42 sp16_42 11.551961
Rsn15_42 sn15_42 sn16_42 11.551961
Rsp15_43 sp15_43 sp16_43 11.551961
Rsn15_43 sn15_43 sn16_43 11.551961
Rsp15_44 sp15_44 sp16_44 11.551961
Rsn15_44 sn15_44 sn16_44 11.551961
Rsp15_45 sp15_45 sp16_45 11.551961
Rsn15_45 sn15_45 sn16_45 11.551961
Rsp15_46 sp15_46 sp16_46 11.551961
Rsn15_46 sn15_46 sn16_46 11.551961
Rsp15_47 sp15_47 sp16_47 11.551961
Rsn15_47 sn15_47 sn16_47 11.551961
Rsp15_48 sp15_48 sp16_48 11.551961
Rsn15_48 sn15_48 sn16_48 11.551961
Rsp15_49 sp15_49 sp16_49 11.551961
Rsn15_49 sn15_49 sn16_49 11.551961
Rsp15_50 sp15_50 sp16_50 11.551961
Rsn15_50 sn15_50 sn16_50 11.551961
Rsp15_51 sp15_51 sp16_51 11.551961
Rsn15_51 sn15_51 sn16_51 11.551961
Rsp15_52 sp15_52 sp16_52 11.551961
Rsn15_52 sn15_52 sn16_52 11.551961
Rsp15_53 sp15_53 sp16_53 11.551961
Rsn15_53 sn15_53 sn16_53 11.551961
Rsp15_54 sp15_54 sp16_54 11.551961
Rsn15_54 sn15_54 sn16_54 11.551961
Rsp15_55 sp15_55 sp16_55 11.551961
Rsn15_55 sn15_55 sn16_55 11.551961
Rsp15_56 sp15_56 sp16_56 11.551961
Rsn15_56 sn15_56 sn16_56 11.551961
Rsp15_57 sp15_57 sp16_57 11.551961
Rsn15_57 sn15_57 sn16_57 11.551961
Rsp15_58 sp15_58 sp16_58 11.551961
Rsn15_58 sn15_58 sn16_58 11.551961
Rsp15_59 sp15_59 sp16_59 11.551961
Rsn15_59 sn15_59 sn16_59 11.551961
Rsp15_60 sp15_60 sp16_60 11.551961
Rsn15_60 sn15_60 sn16_60 11.551961
Rsp15_61 sp15_61 sp16_61 11.551961
Rsn15_61 sn15_61 sn16_61 11.551961
Rsp15_62 sp15_62 sp16_62 11.551961
Rsn15_62 sn15_62 sn16_62 11.551961
Rsp15_63 sp15_63 sp16_63 11.551961
Rsn15_63 sn15_63 sn16_63 11.551961
Rsp15_64 sp15_64 sp16_64 11.551961
Rsn15_64 sn15_64 sn16_64 11.551961
Rsp15_65 sp15_65 sp16_65 11.551961
Rsn15_65 sn15_65 sn16_65 11.551961
Rsp15_66 sp15_66 sp16_66 11.551961
Rsn15_66 sn15_66 sn16_66 11.551961
Rsp15_67 sp15_67 sp16_67 11.551961
Rsn15_67 sn15_67 sn16_67 11.551961
Rsp15_68 sp15_68 sp16_68 11.551961
Rsn15_68 sn15_68 sn16_68 11.551961
Rsp15_69 sp15_69 sp16_69 11.551961
Rsn15_69 sn15_69 sn16_69 11.551961
Rsp15_70 sp15_70 sp16_70 11.551961
Rsn15_70 sn15_70 sn16_70 11.551961
Rsp15_71 sp15_71 sp16_71 11.551961
Rsn15_71 sn15_71 sn16_71 11.551961
Rsp15_72 sp15_72 sp16_72 11.551961
Rsn15_72 sn15_72 sn16_72 11.551961
Rsp15_73 sp15_73 sp16_73 11.551961
Rsn15_73 sn15_73 sn16_73 11.551961
Rsp15_74 sp15_74 sp16_74 11.551961
Rsn15_74 sn15_74 sn16_74 11.551961
Rsp15_75 sp15_75 sp16_75 11.551961
Rsn15_75 sn15_75 sn16_75 11.551961
Rsp15_76 sp15_76 sp16_76 11.551961
Rsn15_76 sn15_76 sn16_76 11.551961
Rsp15_77 sp15_77 sp16_77 11.551961
Rsn15_77 sn15_77 sn16_77 11.551961
Rsp15_78 sp15_78 sp16_78 11.551961
Rsn15_78 sn15_78 sn16_78 11.551961
Rsp15_79 sp15_79 sp16_79 11.551961
Rsn15_79 sn15_79 sn16_79 11.551961
Rsp15_80 sp15_80 sp16_80 11.551961
Rsn15_80 sn15_80 sn16_80 11.551961
Rsp15_81 sp15_81 sp16_81 11.551961
Rsn15_81 sn15_81 sn16_81 11.551961
Rsp15_82 sp15_82 sp16_82 11.551961
Rsn15_82 sn15_82 sn16_82 11.551961
Rsp15_83 sp15_83 sp16_83 11.551961
Rsn15_83 sn15_83 sn16_83 11.551961
Rsp15_84 sp15_84 sp16_84 11.551961
Rsn15_84 sn15_84 sn16_84 11.551961
Rsp16_1 sp16_1 sp17_1 11.551961
Rsn16_1 sn16_1 sn17_1 11.551961
Rsp16_2 sp16_2 sp17_2 11.551961
Rsn16_2 sn16_2 sn17_2 11.551961
Rsp16_3 sp16_3 sp17_3 11.551961
Rsn16_3 sn16_3 sn17_3 11.551961
Rsp16_4 sp16_4 sp17_4 11.551961
Rsn16_4 sn16_4 sn17_4 11.551961
Rsp16_5 sp16_5 sp17_5 11.551961
Rsn16_5 sn16_5 sn17_5 11.551961
Rsp16_6 sp16_6 sp17_6 11.551961
Rsn16_6 sn16_6 sn17_6 11.551961
Rsp16_7 sp16_7 sp17_7 11.551961
Rsn16_7 sn16_7 sn17_7 11.551961
Rsp16_8 sp16_8 sp17_8 11.551961
Rsn16_8 sn16_8 sn17_8 11.551961
Rsp16_9 sp16_9 sp17_9 11.551961
Rsn16_9 sn16_9 sn17_9 11.551961
Rsp16_10 sp16_10 sp17_10 11.551961
Rsn16_10 sn16_10 sn17_10 11.551961
Rsp16_11 sp16_11 sp17_11 11.551961
Rsn16_11 sn16_11 sn17_11 11.551961
Rsp16_12 sp16_12 sp17_12 11.551961
Rsn16_12 sn16_12 sn17_12 11.551961
Rsp16_13 sp16_13 sp17_13 11.551961
Rsn16_13 sn16_13 sn17_13 11.551961
Rsp16_14 sp16_14 sp17_14 11.551961
Rsn16_14 sn16_14 sn17_14 11.551961
Rsp16_15 sp16_15 sp17_15 11.551961
Rsn16_15 sn16_15 sn17_15 11.551961
Rsp16_16 sp16_16 sp17_16 11.551961
Rsn16_16 sn16_16 sn17_16 11.551961
Rsp16_17 sp16_17 sp17_17 11.551961
Rsn16_17 sn16_17 sn17_17 11.551961
Rsp16_18 sp16_18 sp17_18 11.551961
Rsn16_18 sn16_18 sn17_18 11.551961
Rsp16_19 sp16_19 sp17_19 11.551961
Rsn16_19 sn16_19 sn17_19 11.551961
Rsp16_20 sp16_20 sp17_20 11.551961
Rsn16_20 sn16_20 sn17_20 11.551961
Rsp16_21 sp16_21 sp17_21 11.551961
Rsn16_21 sn16_21 sn17_21 11.551961
Rsp16_22 sp16_22 sp17_22 11.551961
Rsn16_22 sn16_22 sn17_22 11.551961
Rsp16_23 sp16_23 sp17_23 11.551961
Rsn16_23 sn16_23 sn17_23 11.551961
Rsp16_24 sp16_24 sp17_24 11.551961
Rsn16_24 sn16_24 sn17_24 11.551961
Rsp16_25 sp16_25 sp17_25 11.551961
Rsn16_25 sn16_25 sn17_25 11.551961
Rsp16_26 sp16_26 sp17_26 11.551961
Rsn16_26 sn16_26 sn17_26 11.551961
Rsp16_27 sp16_27 sp17_27 11.551961
Rsn16_27 sn16_27 sn17_27 11.551961
Rsp16_28 sp16_28 sp17_28 11.551961
Rsn16_28 sn16_28 sn17_28 11.551961
Rsp16_29 sp16_29 sp17_29 11.551961
Rsn16_29 sn16_29 sn17_29 11.551961
Rsp16_30 sp16_30 sp17_30 11.551961
Rsn16_30 sn16_30 sn17_30 11.551961
Rsp16_31 sp16_31 sp17_31 11.551961
Rsn16_31 sn16_31 sn17_31 11.551961
Rsp16_32 sp16_32 sp17_32 11.551961
Rsn16_32 sn16_32 sn17_32 11.551961
Rsp16_33 sp16_33 sp17_33 11.551961
Rsn16_33 sn16_33 sn17_33 11.551961
Rsp16_34 sp16_34 sp17_34 11.551961
Rsn16_34 sn16_34 sn17_34 11.551961
Rsp16_35 sp16_35 sp17_35 11.551961
Rsn16_35 sn16_35 sn17_35 11.551961
Rsp16_36 sp16_36 sp17_36 11.551961
Rsn16_36 sn16_36 sn17_36 11.551961
Rsp16_37 sp16_37 sp17_37 11.551961
Rsn16_37 sn16_37 sn17_37 11.551961
Rsp16_38 sp16_38 sp17_38 11.551961
Rsn16_38 sn16_38 sn17_38 11.551961
Rsp16_39 sp16_39 sp17_39 11.551961
Rsn16_39 sn16_39 sn17_39 11.551961
Rsp16_40 sp16_40 sp17_40 11.551961
Rsn16_40 sn16_40 sn17_40 11.551961
Rsp16_41 sp16_41 sp17_41 11.551961
Rsn16_41 sn16_41 sn17_41 11.551961
Rsp16_42 sp16_42 sp17_42 11.551961
Rsn16_42 sn16_42 sn17_42 11.551961
Rsp16_43 sp16_43 sp17_43 11.551961
Rsn16_43 sn16_43 sn17_43 11.551961
Rsp16_44 sp16_44 sp17_44 11.551961
Rsn16_44 sn16_44 sn17_44 11.551961
Rsp16_45 sp16_45 sp17_45 11.551961
Rsn16_45 sn16_45 sn17_45 11.551961
Rsp16_46 sp16_46 sp17_46 11.551961
Rsn16_46 sn16_46 sn17_46 11.551961
Rsp16_47 sp16_47 sp17_47 11.551961
Rsn16_47 sn16_47 sn17_47 11.551961
Rsp16_48 sp16_48 sp17_48 11.551961
Rsn16_48 sn16_48 sn17_48 11.551961
Rsp16_49 sp16_49 sp17_49 11.551961
Rsn16_49 sn16_49 sn17_49 11.551961
Rsp16_50 sp16_50 sp17_50 11.551961
Rsn16_50 sn16_50 sn17_50 11.551961
Rsp16_51 sp16_51 sp17_51 11.551961
Rsn16_51 sn16_51 sn17_51 11.551961
Rsp16_52 sp16_52 sp17_52 11.551961
Rsn16_52 sn16_52 sn17_52 11.551961
Rsp16_53 sp16_53 sp17_53 11.551961
Rsn16_53 sn16_53 sn17_53 11.551961
Rsp16_54 sp16_54 sp17_54 11.551961
Rsn16_54 sn16_54 sn17_54 11.551961
Rsp16_55 sp16_55 sp17_55 11.551961
Rsn16_55 sn16_55 sn17_55 11.551961
Rsp16_56 sp16_56 sp17_56 11.551961
Rsn16_56 sn16_56 sn17_56 11.551961
Rsp16_57 sp16_57 sp17_57 11.551961
Rsn16_57 sn16_57 sn17_57 11.551961
Rsp16_58 sp16_58 sp17_58 11.551961
Rsn16_58 sn16_58 sn17_58 11.551961
Rsp16_59 sp16_59 sp17_59 11.551961
Rsn16_59 sn16_59 sn17_59 11.551961
Rsp16_60 sp16_60 sp17_60 11.551961
Rsn16_60 sn16_60 sn17_60 11.551961
Rsp16_61 sp16_61 sp17_61 11.551961
Rsn16_61 sn16_61 sn17_61 11.551961
Rsp16_62 sp16_62 sp17_62 11.551961
Rsn16_62 sn16_62 sn17_62 11.551961
Rsp16_63 sp16_63 sp17_63 11.551961
Rsn16_63 sn16_63 sn17_63 11.551961
Rsp16_64 sp16_64 sp17_64 11.551961
Rsn16_64 sn16_64 sn17_64 11.551961
Rsp16_65 sp16_65 sp17_65 11.551961
Rsn16_65 sn16_65 sn17_65 11.551961
Rsp16_66 sp16_66 sp17_66 11.551961
Rsn16_66 sn16_66 sn17_66 11.551961
Rsp16_67 sp16_67 sp17_67 11.551961
Rsn16_67 sn16_67 sn17_67 11.551961
Rsp16_68 sp16_68 sp17_68 11.551961
Rsn16_68 sn16_68 sn17_68 11.551961
Rsp16_69 sp16_69 sp17_69 11.551961
Rsn16_69 sn16_69 sn17_69 11.551961
Rsp16_70 sp16_70 sp17_70 11.551961
Rsn16_70 sn16_70 sn17_70 11.551961
Rsp16_71 sp16_71 sp17_71 11.551961
Rsn16_71 sn16_71 sn17_71 11.551961
Rsp16_72 sp16_72 sp17_72 11.551961
Rsn16_72 sn16_72 sn17_72 11.551961
Rsp16_73 sp16_73 sp17_73 11.551961
Rsn16_73 sn16_73 sn17_73 11.551961
Rsp16_74 sp16_74 sp17_74 11.551961
Rsn16_74 sn16_74 sn17_74 11.551961
Rsp16_75 sp16_75 sp17_75 11.551961
Rsn16_75 sn16_75 sn17_75 11.551961
Rsp16_76 sp16_76 sp17_76 11.551961
Rsn16_76 sn16_76 sn17_76 11.551961
Rsp16_77 sp16_77 sp17_77 11.551961
Rsn16_77 sn16_77 sn17_77 11.551961
Rsp16_78 sp16_78 sp17_78 11.551961
Rsn16_78 sn16_78 sn17_78 11.551961
Rsp16_79 sp16_79 sp17_79 11.551961
Rsn16_79 sn16_79 sn17_79 11.551961
Rsp16_80 sp16_80 sp17_80 11.551961
Rsn16_80 sn16_80 sn17_80 11.551961
Rsp16_81 sp16_81 sp17_81 11.551961
Rsn16_81 sn16_81 sn17_81 11.551961
Rsp16_82 sp16_82 sp17_82 11.551961
Rsn16_82 sn16_82 sn17_82 11.551961
Rsp16_83 sp16_83 sp17_83 11.551961
Rsn16_83 sn16_83 sn17_83 11.551961
Rsp16_84 sp16_84 sp17_84 11.551961
Rsn16_84 sn16_84 sn17_84 11.551961
Rsp17_1 sp17_1 sp18_1 11.551961
Rsn17_1 sn17_1 sn18_1 11.551961
Rsp17_2 sp17_2 sp18_2 11.551961
Rsn17_2 sn17_2 sn18_2 11.551961
Rsp17_3 sp17_3 sp18_3 11.551961
Rsn17_3 sn17_3 sn18_3 11.551961
Rsp17_4 sp17_4 sp18_4 11.551961
Rsn17_4 sn17_4 sn18_4 11.551961
Rsp17_5 sp17_5 sp18_5 11.551961
Rsn17_5 sn17_5 sn18_5 11.551961
Rsp17_6 sp17_6 sp18_6 11.551961
Rsn17_6 sn17_6 sn18_6 11.551961
Rsp17_7 sp17_7 sp18_7 11.551961
Rsn17_7 sn17_7 sn18_7 11.551961
Rsp17_8 sp17_8 sp18_8 11.551961
Rsn17_8 sn17_8 sn18_8 11.551961
Rsp17_9 sp17_9 sp18_9 11.551961
Rsn17_9 sn17_9 sn18_9 11.551961
Rsp17_10 sp17_10 sp18_10 11.551961
Rsn17_10 sn17_10 sn18_10 11.551961
Rsp17_11 sp17_11 sp18_11 11.551961
Rsn17_11 sn17_11 sn18_11 11.551961
Rsp17_12 sp17_12 sp18_12 11.551961
Rsn17_12 sn17_12 sn18_12 11.551961
Rsp17_13 sp17_13 sp18_13 11.551961
Rsn17_13 sn17_13 sn18_13 11.551961
Rsp17_14 sp17_14 sp18_14 11.551961
Rsn17_14 sn17_14 sn18_14 11.551961
Rsp17_15 sp17_15 sp18_15 11.551961
Rsn17_15 sn17_15 sn18_15 11.551961
Rsp17_16 sp17_16 sp18_16 11.551961
Rsn17_16 sn17_16 sn18_16 11.551961
Rsp17_17 sp17_17 sp18_17 11.551961
Rsn17_17 sn17_17 sn18_17 11.551961
Rsp17_18 sp17_18 sp18_18 11.551961
Rsn17_18 sn17_18 sn18_18 11.551961
Rsp17_19 sp17_19 sp18_19 11.551961
Rsn17_19 sn17_19 sn18_19 11.551961
Rsp17_20 sp17_20 sp18_20 11.551961
Rsn17_20 sn17_20 sn18_20 11.551961
Rsp17_21 sp17_21 sp18_21 11.551961
Rsn17_21 sn17_21 sn18_21 11.551961
Rsp17_22 sp17_22 sp18_22 11.551961
Rsn17_22 sn17_22 sn18_22 11.551961
Rsp17_23 sp17_23 sp18_23 11.551961
Rsn17_23 sn17_23 sn18_23 11.551961
Rsp17_24 sp17_24 sp18_24 11.551961
Rsn17_24 sn17_24 sn18_24 11.551961
Rsp17_25 sp17_25 sp18_25 11.551961
Rsn17_25 sn17_25 sn18_25 11.551961
Rsp17_26 sp17_26 sp18_26 11.551961
Rsn17_26 sn17_26 sn18_26 11.551961
Rsp17_27 sp17_27 sp18_27 11.551961
Rsn17_27 sn17_27 sn18_27 11.551961
Rsp17_28 sp17_28 sp18_28 11.551961
Rsn17_28 sn17_28 sn18_28 11.551961
Rsp17_29 sp17_29 sp18_29 11.551961
Rsn17_29 sn17_29 sn18_29 11.551961
Rsp17_30 sp17_30 sp18_30 11.551961
Rsn17_30 sn17_30 sn18_30 11.551961
Rsp17_31 sp17_31 sp18_31 11.551961
Rsn17_31 sn17_31 sn18_31 11.551961
Rsp17_32 sp17_32 sp18_32 11.551961
Rsn17_32 sn17_32 sn18_32 11.551961
Rsp17_33 sp17_33 sp18_33 11.551961
Rsn17_33 sn17_33 sn18_33 11.551961
Rsp17_34 sp17_34 sp18_34 11.551961
Rsn17_34 sn17_34 sn18_34 11.551961
Rsp17_35 sp17_35 sp18_35 11.551961
Rsn17_35 sn17_35 sn18_35 11.551961
Rsp17_36 sp17_36 sp18_36 11.551961
Rsn17_36 sn17_36 sn18_36 11.551961
Rsp17_37 sp17_37 sp18_37 11.551961
Rsn17_37 sn17_37 sn18_37 11.551961
Rsp17_38 sp17_38 sp18_38 11.551961
Rsn17_38 sn17_38 sn18_38 11.551961
Rsp17_39 sp17_39 sp18_39 11.551961
Rsn17_39 sn17_39 sn18_39 11.551961
Rsp17_40 sp17_40 sp18_40 11.551961
Rsn17_40 sn17_40 sn18_40 11.551961
Rsp17_41 sp17_41 sp18_41 11.551961
Rsn17_41 sn17_41 sn18_41 11.551961
Rsp17_42 sp17_42 sp18_42 11.551961
Rsn17_42 sn17_42 sn18_42 11.551961
Rsp17_43 sp17_43 sp18_43 11.551961
Rsn17_43 sn17_43 sn18_43 11.551961
Rsp17_44 sp17_44 sp18_44 11.551961
Rsn17_44 sn17_44 sn18_44 11.551961
Rsp17_45 sp17_45 sp18_45 11.551961
Rsn17_45 sn17_45 sn18_45 11.551961
Rsp17_46 sp17_46 sp18_46 11.551961
Rsn17_46 sn17_46 sn18_46 11.551961
Rsp17_47 sp17_47 sp18_47 11.551961
Rsn17_47 sn17_47 sn18_47 11.551961
Rsp17_48 sp17_48 sp18_48 11.551961
Rsn17_48 sn17_48 sn18_48 11.551961
Rsp17_49 sp17_49 sp18_49 11.551961
Rsn17_49 sn17_49 sn18_49 11.551961
Rsp17_50 sp17_50 sp18_50 11.551961
Rsn17_50 sn17_50 sn18_50 11.551961
Rsp17_51 sp17_51 sp18_51 11.551961
Rsn17_51 sn17_51 sn18_51 11.551961
Rsp17_52 sp17_52 sp18_52 11.551961
Rsn17_52 sn17_52 sn18_52 11.551961
Rsp17_53 sp17_53 sp18_53 11.551961
Rsn17_53 sn17_53 sn18_53 11.551961
Rsp17_54 sp17_54 sp18_54 11.551961
Rsn17_54 sn17_54 sn18_54 11.551961
Rsp17_55 sp17_55 sp18_55 11.551961
Rsn17_55 sn17_55 sn18_55 11.551961
Rsp17_56 sp17_56 sp18_56 11.551961
Rsn17_56 sn17_56 sn18_56 11.551961
Rsp17_57 sp17_57 sp18_57 11.551961
Rsn17_57 sn17_57 sn18_57 11.551961
Rsp17_58 sp17_58 sp18_58 11.551961
Rsn17_58 sn17_58 sn18_58 11.551961
Rsp17_59 sp17_59 sp18_59 11.551961
Rsn17_59 sn17_59 sn18_59 11.551961
Rsp17_60 sp17_60 sp18_60 11.551961
Rsn17_60 sn17_60 sn18_60 11.551961
Rsp17_61 sp17_61 sp18_61 11.551961
Rsn17_61 sn17_61 sn18_61 11.551961
Rsp17_62 sp17_62 sp18_62 11.551961
Rsn17_62 sn17_62 sn18_62 11.551961
Rsp17_63 sp17_63 sp18_63 11.551961
Rsn17_63 sn17_63 sn18_63 11.551961
Rsp17_64 sp17_64 sp18_64 11.551961
Rsn17_64 sn17_64 sn18_64 11.551961
Rsp17_65 sp17_65 sp18_65 11.551961
Rsn17_65 sn17_65 sn18_65 11.551961
Rsp17_66 sp17_66 sp18_66 11.551961
Rsn17_66 sn17_66 sn18_66 11.551961
Rsp17_67 sp17_67 sp18_67 11.551961
Rsn17_67 sn17_67 sn18_67 11.551961
Rsp17_68 sp17_68 sp18_68 11.551961
Rsn17_68 sn17_68 sn18_68 11.551961
Rsp17_69 sp17_69 sp18_69 11.551961
Rsn17_69 sn17_69 sn18_69 11.551961
Rsp17_70 sp17_70 sp18_70 11.551961
Rsn17_70 sn17_70 sn18_70 11.551961
Rsp17_71 sp17_71 sp18_71 11.551961
Rsn17_71 sn17_71 sn18_71 11.551961
Rsp17_72 sp17_72 sp18_72 11.551961
Rsn17_72 sn17_72 sn18_72 11.551961
Rsp17_73 sp17_73 sp18_73 11.551961
Rsn17_73 sn17_73 sn18_73 11.551961
Rsp17_74 sp17_74 sp18_74 11.551961
Rsn17_74 sn17_74 sn18_74 11.551961
Rsp17_75 sp17_75 sp18_75 11.551961
Rsn17_75 sn17_75 sn18_75 11.551961
Rsp17_76 sp17_76 sp18_76 11.551961
Rsn17_76 sn17_76 sn18_76 11.551961
Rsp17_77 sp17_77 sp18_77 11.551961
Rsn17_77 sn17_77 sn18_77 11.551961
Rsp17_78 sp17_78 sp18_78 11.551961
Rsn17_78 sn17_78 sn18_78 11.551961
Rsp17_79 sp17_79 sp18_79 11.551961
Rsn17_79 sn17_79 sn18_79 11.551961
Rsp17_80 sp17_80 sp18_80 11.551961
Rsn17_80 sn17_80 sn18_80 11.551961
Rsp17_81 sp17_81 sp18_81 11.551961
Rsn17_81 sn17_81 sn18_81 11.551961
Rsp17_82 sp17_82 sp18_82 11.551961
Rsn17_82 sn17_82 sn18_82 11.551961
Rsp17_83 sp17_83 sp18_83 11.551961
Rsn17_83 sn17_83 sn18_83 11.551961
Rsp17_84 sp17_84 sp18_84 11.551961
Rsn17_84 sn17_84 sn18_84 11.551961
Rsp18_1 sp18_1 sp19_1 11.551961
Rsn18_1 sn18_1 sn19_1 11.551961
Rsp18_2 sp18_2 sp19_2 11.551961
Rsn18_2 sn18_2 sn19_2 11.551961
Rsp18_3 sp18_3 sp19_3 11.551961
Rsn18_3 sn18_3 sn19_3 11.551961
Rsp18_4 sp18_4 sp19_4 11.551961
Rsn18_4 sn18_4 sn19_4 11.551961
Rsp18_5 sp18_5 sp19_5 11.551961
Rsn18_5 sn18_5 sn19_5 11.551961
Rsp18_6 sp18_6 sp19_6 11.551961
Rsn18_6 sn18_6 sn19_6 11.551961
Rsp18_7 sp18_7 sp19_7 11.551961
Rsn18_7 sn18_7 sn19_7 11.551961
Rsp18_8 sp18_8 sp19_8 11.551961
Rsn18_8 sn18_8 sn19_8 11.551961
Rsp18_9 sp18_9 sp19_9 11.551961
Rsn18_9 sn18_9 sn19_9 11.551961
Rsp18_10 sp18_10 sp19_10 11.551961
Rsn18_10 sn18_10 sn19_10 11.551961
Rsp18_11 sp18_11 sp19_11 11.551961
Rsn18_11 sn18_11 sn19_11 11.551961
Rsp18_12 sp18_12 sp19_12 11.551961
Rsn18_12 sn18_12 sn19_12 11.551961
Rsp18_13 sp18_13 sp19_13 11.551961
Rsn18_13 sn18_13 sn19_13 11.551961
Rsp18_14 sp18_14 sp19_14 11.551961
Rsn18_14 sn18_14 sn19_14 11.551961
Rsp18_15 sp18_15 sp19_15 11.551961
Rsn18_15 sn18_15 sn19_15 11.551961
Rsp18_16 sp18_16 sp19_16 11.551961
Rsn18_16 sn18_16 sn19_16 11.551961
Rsp18_17 sp18_17 sp19_17 11.551961
Rsn18_17 sn18_17 sn19_17 11.551961
Rsp18_18 sp18_18 sp19_18 11.551961
Rsn18_18 sn18_18 sn19_18 11.551961
Rsp18_19 sp18_19 sp19_19 11.551961
Rsn18_19 sn18_19 sn19_19 11.551961
Rsp18_20 sp18_20 sp19_20 11.551961
Rsn18_20 sn18_20 sn19_20 11.551961
Rsp18_21 sp18_21 sp19_21 11.551961
Rsn18_21 sn18_21 sn19_21 11.551961
Rsp18_22 sp18_22 sp19_22 11.551961
Rsn18_22 sn18_22 sn19_22 11.551961
Rsp18_23 sp18_23 sp19_23 11.551961
Rsn18_23 sn18_23 sn19_23 11.551961
Rsp18_24 sp18_24 sp19_24 11.551961
Rsn18_24 sn18_24 sn19_24 11.551961
Rsp18_25 sp18_25 sp19_25 11.551961
Rsn18_25 sn18_25 sn19_25 11.551961
Rsp18_26 sp18_26 sp19_26 11.551961
Rsn18_26 sn18_26 sn19_26 11.551961
Rsp18_27 sp18_27 sp19_27 11.551961
Rsn18_27 sn18_27 sn19_27 11.551961
Rsp18_28 sp18_28 sp19_28 11.551961
Rsn18_28 sn18_28 sn19_28 11.551961
Rsp18_29 sp18_29 sp19_29 11.551961
Rsn18_29 sn18_29 sn19_29 11.551961
Rsp18_30 sp18_30 sp19_30 11.551961
Rsn18_30 sn18_30 sn19_30 11.551961
Rsp18_31 sp18_31 sp19_31 11.551961
Rsn18_31 sn18_31 sn19_31 11.551961
Rsp18_32 sp18_32 sp19_32 11.551961
Rsn18_32 sn18_32 sn19_32 11.551961
Rsp18_33 sp18_33 sp19_33 11.551961
Rsn18_33 sn18_33 sn19_33 11.551961
Rsp18_34 sp18_34 sp19_34 11.551961
Rsn18_34 sn18_34 sn19_34 11.551961
Rsp18_35 sp18_35 sp19_35 11.551961
Rsn18_35 sn18_35 sn19_35 11.551961
Rsp18_36 sp18_36 sp19_36 11.551961
Rsn18_36 sn18_36 sn19_36 11.551961
Rsp18_37 sp18_37 sp19_37 11.551961
Rsn18_37 sn18_37 sn19_37 11.551961
Rsp18_38 sp18_38 sp19_38 11.551961
Rsn18_38 sn18_38 sn19_38 11.551961
Rsp18_39 sp18_39 sp19_39 11.551961
Rsn18_39 sn18_39 sn19_39 11.551961
Rsp18_40 sp18_40 sp19_40 11.551961
Rsn18_40 sn18_40 sn19_40 11.551961
Rsp18_41 sp18_41 sp19_41 11.551961
Rsn18_41 sn18_41 sn19_41 11.551961
Rsp18_42 sp18_42 sp19_42 11.551961
Rsn18_42 sn18_42 sn19_42 11.551961
Rsp18_43 sp18_43 sp19_43 11.551961
Rsn18_43 sn18_43 sn19_43 11.551961
Rsp18_44 sp18_44 sp19_44 11.551961
Rsn18_44 sn18_44 sn19_44 11.551961
Rsp18_45 sp18_45 sp19_45 11.551961
Rsn18_45 sn18_45 sn19_45 11.551961
Rsp18_46 sp18_46 sp19_46 11.551961
Rsn18_46 sn18_46 sn19_46 11.551961
Rsp18_47 sp18_47 sp19_47 11.551961
Rsn18_47 sn18_47 sn19_47 11.551961
Rsp18_48 sp18_48 sp19_48 11.551961
Rsn18_48 sn18_48 sn19_48 11.551961
Rsp18_49 sp18_49 sp19_49 11.551961
Rsn18_49 sn18_49 sn19_49 11.551961
Rsp18_50 sp18_50 sp19_50 11.551961
Rsn18_50 sn18_50 sn19_50 11.551961
Rsp18_51 sp18_51 sp19_51 11.551961
Rsn18_51 sn18_51 sn19_51 11.551961
Rsp18_52 sp18_52 sp19_52 11.551961
Rsn18_52 sn18_52 sn19_52 11.551961
Rsp18_53 sp18_53 sp19_53 11.551961
Rsn18_53 sn18_53 sn19_53 11.551961
Rsp18_54 sp18_54 sp19_54 11.551961
Rsn18_54 sn18_54 sn19_54 11.551961
Rsp18_55 sp18_55 sp19_55 11.551961
Rsn18_55 sn18_55 sn19_55 11.551961
Rsp18_56 sp18_56 sp19_56 11.551961
Rsn18_56 sn18_56 sn19_56 11.551961
Rsp18_57 sp18_57 sp19_57 11.551961
Rsn18_57 sn18_57 sn19_57 11.551961
Rsp18_58 sp18_58 sp19_58 11.551961
Rsn18_58 sn18_58 sn19_58 11.551961
Rsp18_59 sp18_59 sp19_59 11.551961
Rsn18_59 sn18_59 sn19_59 11.551961
Rsp18_60 sp18_60 sp19_60 11.551961
Rsn18_60 sn18_60 sn19_60 11.551961
Rsp18_61 sp18_61 sp19_61 11.551961
Rsn18_61 sn18_61 sn19_61 11.551961
Rsp18_62 sp18_62 sp19_62 11.551961
Rsn18_62 sn18_62 sn19_62 11.551961
Rsp18_63 sp18_63 sp19_63 11.551961
Rsn18_63 sn18_63 sn19_63 11.551961
Rsp18_64 sp18_64 sp19_64 11.551961
Rsn18_64 sn18_64 sn19_64 11.551961
Rsp18_65 sp18_65 sp19_65 11.551961
Rsn18_65 sn18_65 sn19_65 11.551961
Rsp18_66 sp18_66 sp19_66 11.551961
Rsn18_66 sn18_66 sn19_66 11.551961
Rsp18_67 sp18_67 sp19_67 11.551961
Rsn18_67 sn18_67 sn19_67 11.551961
Rsp18_68 sp18_68 sp19_68 11.551961
Rsn18_68 sn18_68 sn19_68 11.551961
Rsp18_69 sp18_69 sp19_69 11.551961
Rsn18_69 sn18_69 sn19_69 11.551961
Rsp18_70 sp18_70 sp19_70 11.551961
Rsn18_70 sn18_70 sn19_70 11.551961
Rsp18_71 sp18_71 sp19_71 11.551961
Rsn18_71 sn18_71 sn19_71 11.551961
Rsp18_72 sp18_72 sp19_72 11.551961
Rsn18_72 sn18_72 sn19_72 11.551961
Rsp18_73 sp18_73 sp19_73 11.551961
Rsn18_73 sn18_73 sn19_73 11.551961
Rsp18_74 sp18_74 sp19_74 11.551961
Rsn18_74 sn18_74 sn19_74 11.551961
Rsp18_75 sp18_75 sp19_75 11.551961
Rsn18_75 sn18_75 sn19_75 11.551961
Rsp18_76 sp18_76 sp19_76 11.551961
Rsn18_76 sn18_76 sn19_76 11.551961
Rsp18_77 sp18_77 sp19_77 11.551961
Rsn18_77 sn18_77 sn19_77 11.551961
Rsp18_78 sp18_78 sp19_78 11.551961
Rsn18_78 sn18_78 sn19_78 11.551961
Rsp18_79 sp18_79 sp19_79 11.551961
Rsn18_79 sn18_79 sn19_79 11.551961
Rsp18_80 sp18_80 sp19_80 11.551961
Rsn18_80 sn18_80 sn19_80 11.551961
Rsp18_81 sp18_81 sp19_81 11.551961
Rsn18_81 sn18_81 sn19_81 11.551961
Rsp18_82 sp18_82 sp19_82 11.551961
Rsn18_82 sn18_82 sn19_82 11.551961
Rsp18_83 sp18_83 sp19_83 11.551961
Rsn18_83 sn18_83 sn19_83 11.551961
Rsp18_84 sp18_84 sp19_84 11.551961
Rsn18_84 sn18_84 sn19_84 11.551961
Rsp19_1 sp19_1 sp20_1 11.551961
Rsn19_1 sn19_1 sn20_1 11.551961
Rsp19_2 sp19_2 sp20_2 11.551961
Rsn19_2 sn19_2 sn20_2 11.551961
Rsp19_3 sp19_3 sp20_3 11.551961
Rsn19_3 sn19_3 sn20_3 11.551961
Rsp19_4 sp19_4 sp20_4 11.551961
Rsn19_4 sn19_4 sn20_4 11.551961
Rsp19_5 sp19_5 sp20_5 11.551961
Rsn19_5 sn19_5 sn20_5 11.551961
Rsp19_6 sp19_6 sp20_6 11.551961
Rsn19_6 sn19_6 sn20_6 11.551961
Rsp19_7 sp19_7 sp20_7 11.551961
Rsn19_7 sn19_7 sn20_7 11.551961
Rsp19_8 sp19_8 sp20_8 11.551961
Rsn19_8 sn19_8 sn20_8 11.551961
Rsp19_9 sp19_9 sp20_9 11.551961
Rsn19_9 sn19_9 sn20_9 11.551961
Rsp19_10 sp19_10 sp20_10 11.551961
Rsn19_10 sn19_10 sn20_10 11.551961
Rsp19_11 sp19_11 sp20_11 11.551961
Rsn19_11 sn19_11 sn20_11 11.551961
Rsp19_12 sp19_12 sp20_12 11.551961
Rsn19_12 sn19_12 sn20_12 11.551961
Rsp19_13 sp19_13 sp20_13 11.551961
Rsn19_13 sn19_13 sn20_13 11.551961
Rsp19_14 sp19_14 sp20_14 11.551961
Rsn19_14 sn19_14 sn20_14 11.551961
Rsp19_15 sp19_15 sp20_15 11.551961
Rsn19_15 sn19_15 sn20_15 11.551961
Rsp19_16 sp19_16 sp20_16 11.551961
Rsn19_16 sn19_16 sn20_16 11.551961
Rsp19_17 sp19_17 sp20_17 11.551961
Rsn19_17 sn19_17 sn20_17 11.551961
Rsp19_18 sp19_18 sp20_18 11.551961
Rsn19_18 sn19_18 sn20_18 11.551961
Rsp19_19 sp19_19 sp20_19 11.551961
Rsn19_19 sn19_19 sn20_19 11.551961
Rsp19_20 sp19_20 sp20_20 11.551961
Rsn19_20 sn19_20 sn20_20 11.551961
Rsp19_21 sp19_21 sp20_21 11.551961
Rsn19_21 sn19_21 sn20_21 11.551961
Rsp19_22 sp19_22 sp20_22 11.551961
Rsn19_22 sn19_22 sn20_22 11.551961
Rsp19_23 sp19_23 sp20_23 11.551961
Rsn19_23 sn19_23 sn20_23 11.551961
Rsp19_24 sp19_24 sp20_24 11.551961
Rsn19_24 sn19_24 sn20_24 11.551961
Rsp19_25 sp19_25 sp20_25 11.551961
Rsn19_25 sn19_25 sn20_25 11.551961
Rsp19_26 sp19_26 sp20_26 11.551961
Rsn19_26 sn19_26 sn20_26 11.551961
Rsp19_27 sp19_27 sp20_27 11.551961
Rsn19_27 sn19_27 sn20_27 11.551961
Rsp19_28 sp19_28 sp20_28 11.551961
Rsn19_28 sn19_28 sn20_28 11.551961
Rsp19_29 sp19_29 sp20_29 11.551961
Rsn19_29 sn19_29 sn20_29 11.551961
Rsp19_30 sp19_30 sp20_30 11.551961
Rsn19_30 sn19_30 sn20_30 11.551961
Rsp19_31 sp19_31 sp20_31 11.551961
Rsn19_31 sn19_31 sn20_31 11.551961
Rsp19_32 sp19_32 sp20_32 11.551961
Rsn19_32 sn19_32 sn20_32 11.551961
Rsp19_33 sp19_33 sp20_33 11.551961
Rsn19_33 sn19_33 sn20_33 11.551961
Rsp19_34 sp19_34 sp20_34 11.551961
Rsn19_34 sn19_34 sn20_34 11.551961
Rsp19_35 sp19_35 sp20_35 11.551961
Rsn19_35 sn19_35 sn20_35 11.551961
Rsp19_36 sp19_36 sp20_36 11.551961
Rsn19_36 sn19_36 sn20_36 11.551961
Rsp19_37 sp19_37 sp20_37 11.551961
Rsn19_37 sn19_37 sn20_37 11.551961
Rsp19_38 sp19_38 sp20_38 11.551961
Rsn19_38 sn19_38 sn20_38 11.551961
Rsp19_39 sp19_39 sp20_39 11.551961
Rsn19_39 sn19_39 sn20_39 11.551961
Rsp19_40 sp19_40 sp20_40 11.551961
Rsn19_40 sn19_40 sn20_40 11.551961
Rsp19_41 sp19_41 sp20_41 11.551961
Rsn19_41 sn19_41 sn20_41 11.551961
Rsp19_42 sp19_42 sp20_42 11.551961
Rsn19_42 sn19_42 sn20_42 11.551961
Rsp19_43 sp19_43 sp20_43 11.551961
Rsn19_43 sn19_43 sn20_43 11.551961
Rsp19_44 sp19_44 sp20_44 11.551961
Rsn19_44 sn19_44 sn20_44 11.551961
Rsp19_45 sp19_45 sp20_45 11.551961
Rsn19_45 sn19_45 sn20_45 11.551961
Rsp19_46 sp19_46 sp20_46 11.551961
Rsn19_46 sn19_46 sn20_46 11.551961
Rsp19_47 sp19_47 sp20_47 11.551961
Rsn19_47 sn19_47 sn20_47 11.551961
Rsp19_48 sp19_48 sp20_48 11.551961
Rsn19_48 sn19_48 sn20_48 11.551961
Rsp19_49 sp19_49 sp20_49 11.551961
Rsn19_49 sn19_49 sn20_49 11.551961
Rsp19_50 sp19_50 sp20_50 11.551961
Rsn19_50 sn19_50 sn20_50 11.551961
Rsp19_51 sp19_51 sp20_51 11.551961
Rsn19_51 sn19_51 sn20_51 11.551961
Rsp19_52 sp19_52 sp20_52 11.551961
Rsn19_52 sn19_52 sn20_52 11.551961
Rsp19_53 sp19_53 sp20_53 11.551961
Rsn19_53 sn19_53 sn20_53 11.551961
Rsp19_54 sp19_54 sp20_54 11.551961
Rsn19_54 sn19_54 sn20_54 11.551961
Rsp19_55 sp19_55 sp20_55 11.551961
Rsn19_55 sn19_55 sn20_55 11.551961
Rsp19_56 sp19_56 sp20_56 11.551961
Rsn19_56 sn19_56 sn20_56 11.551961
Rsp19_57 sp19_57 sp20_57 11.551961
Rsn19_57 sn19_57 sn20_57 11.551961
Rsp19_58 sp19_58 sp20_58 11.551961
Rsn19_58 sn19_58 sn20_58 11.551961
Rsp19_59 sp19_59 sp20_59 11.551961
Rsn19_59 sn19_59 sn20_59 11.551961
Rsp19_60 sp19_60 sp20_60 11.551961
Rsn19_60 sn19_60 sn20_60 11.551961
Rsp19_61 sp19_61 sp20_61 11.551961
Rsn19_61 sn19_61 sn20_61 11.551961
Rsp19_62 sp19_62 sp20_62 11.551961
Rsn19_62 sn19_62 sn20_62 11.551961
Rsp19_63 sp19_63 sp20_63 11.551961
Rsn19_63 sn19_63 sn20_63 11.551961
Rsp19_64 sp19_64 sp20_64 11.551961
Rsn19_64 sn19_64 sn20_64 11.551961
Rsp19_65 sp19_65 sp20_65 11.551961
Rsn19_65 sn19_65 sn20_65 11.551961
Rsp19_66 sp19_66 sp20_66 11.551961
Rsn19_66 sn19_66 sn20_66 11.551961
Rsp19_67 sp19_67 sp20_67 11.551961
Rsn19_67 sn19_67 sn20_67 11.551961
Rsp19_68 sp19_68 sp20_68 11.551961
Rsn19_68 sn19_68 sn20_68 11.551961
Rsp19_69 sp19_69 sp20_69 11.551961
Rsn19_69 sn19_69 sn20_69 11.551961
Rsp19_70 sp19_70 sp20_70 11.551961
Rsn19_70 sn19_70 sn20_70 11.551961
Rsp19_71 sp19_71 sp20_71 11.551961
Rsn19_71 sn19_71 sn20_71 11.551961
Rsp19_72 sp19_72 sp20_72 11.551961
Rsn19_72 sn19_72 sn20_72 11.551961
Rsp19_73 sp19_73 sp20_73 11.551961
Rsn19_73 sn19_73 sn20_73 11.551961
Rsp19_74 sp19_74 sp20_74 11.551961
Rsn19_74 sn19_74 sn20_74 11.551961
Rsp19_75 sp19_75 sp20_75 11.551961
Rsn19_75 sn19_75 sn20_75 11.551961
Rsp19_76 sp19_76 sp20_76 11.551961
Rsn19_76 sn19_76 sn20_76 11.551961
Rsp19_77 sp19_77 sp20_77 11.551961
Rsn19_77 sn19_77 sn20_77 11.551961
Rsp19_78 sp19_78 sp20_78 11.551961
Rsn19_78 sn19_78 sn20_78 11.551961
Rsp19_79 sp19_79 sp20_79 11.551961
Rsn19_79 sn19_79 sn20_79 11.551961
Rsp19_80 sp19_80 sp20_80 11.551961
Rsn19_80 sn19_80 sn20_80 11.551961
Rsp19_81 sp19_81 sp20_81 11.551961
Rsn19_81 sn19_81 sn20_81 11.551961
Rsp19_82 sp19_82 sp20_82 11.551961
Rsn19_82 sn19_82 sn20_82 11.551961
Rsp19_83 sp19_83 sp20_83 11.551961
Rsn19_83 sn19_83 sn20_83 11.551961
Rsp19_84 sp19_84 sp20_84 11.551961
Rsn19_84 sn19_84 sn20_84 11.551961
Rsp20_1 sp20_1 sp21_1 11.551961
Rsn20_1 sn20_1 sn21_1 11.551961
Rsp20_2 sp20_2 sp21_2 11.551961
Rsn20_2 sn20_2 sn21_2 11.551961
Rsp20_3 sp20_3 sp21_3 11.551961
Rsn20_3 sn20_3 sn21_3 11.551961
Rsp20_4 sp20_4 sp21_4 11.551961
Rsn20_4 sn20_4 sn21_4 11.551961
Rsp20_5 sp20_5 sp21_5 11.551961
Rsn20_5 sn20_5 sn21_5 11.551961
Rsp20_6 sp20_6 sp21_6 11.551961
Rsn20_6 sn20_6 sn21_6 11.551961
Rsp20_7 sp20_7 sp21_7 11.551961
Rsn20_7 sn20_7 sn21_7 11.551961
Rsp20_8 sp20_8 sp21_8 11.551961
Rsn20_8 sn20_8 sn21_8 11.551961
Rsp20_9 sp20_9 sp21_9 11.551961
Rsn20_9 sn20_9 sn21_9 11.551961
Rsp20_10 sp20_10 sp21_10 11.551961
Rsn20_10 sn20_10 sn21_10 11.551961
Rsp20_11 sp20_11 sp21_11 11.551961
Rsn20_11 sn20_11 sn21_11 11.551961
Rsp20_12 sp20_12 sp21_12 11.551961
Rsn20_12 sn20_12 sn21_12 11.551961
Rsp20_13 sp20_13 sp21_13 11.551961
Rsn20_13 sn20_13 sn21_13 11.551961
Rsp20_14 sp20_14 sp21_14 11.551961
Rsn20_14 sn20_14 sn21_14 11.551961
Rsp20_15 sp20_15 sp21_15 11.551961
Rsn20_15 sn20_15 sn21_15 11.551961
Rsp20_16 sp20_16 sp21_16 11.551961
Rsn20_16 sn20_16 sn21_16 11.551961
Rsp20_17 sp20_17 sp21_17 11.551961
Rsn20_17 sn20_17 sn21_17 11.551961
Rsp20_18 sp20_18 sp21_18 11.551961
Rsn20_18 sn20_18 sn21_18 11.551961
Rsp20_19 sp20_19 sp21_19 11.551961
Rsn20_19 sn20_19 sn21_19 11.551961
Rsp20_20 sp20_20 sp21_20 11.551961
Rsn20_20 sn20_20 sn21_20 11.551961
Rsp20_21 sp20_21 sp21_21 11.551961
Rsn20_21 sn20_21 sn21_21 11.551961
Rsp20_22 sp20_22 sp21_22 11.551961
Rsn20_22 sn20_22 sn21_22 11.551961
Rsp20_23 sp20_23 sp21_23 11.551961
Rsn20_23 sn20_23 sn21_23 11.551961
Rsp20_24 sp20_24 sp21_24 11.551961
Rsn20_24 sn20_24 sn21_24 11.551961
Rsp20_25 sp20_25 sp21_25 11.551961
Rsn20_25 sn20_25 sn21_25 11.551961
Rsp20_26 sp20_26 sp21_26 11.551961
Rsn20_26 sn20_26 sn21_26 11.551961
Rsp20_27 sp20_27 sp21_27 11.551961
Rsn20_27 sn20_27 sn21_27 11.551961
Rsp20_28 sp20_28 sp21_28 11.551961
Rsn20_28 sn20_28 sn21_28 11.551961
Rsp20_29 sp20_29 sp21_29 11.551961
Rsn20_29 sn20_29 sn21_29 11.551961
Rsp20_30 sp20_30 sp21_30 11.551961
Rsn20_30 sn20_30 sn21_30 11.551961
Rsp20_31 sp20_31 sp21_31 11.551961
Rsn20_31 sn20_31 sn21_31 11.551961
Rsp20_32 sp20_32 sp21_32 11.551961
Rsn20_32 sn20_32 sn21_32 11.551961
Rsp20_33 sp20_33 sp21_33 11.551961
Rsn20_33 sn20_33 sn21_33 11.551961
Rsp20_34 sp20_34 sp21_34 11.551961
Rsn20_34 sn20_34 sn21_34 11.551961
Rsp20_35 sp20_35 sp21_35 11.551961
Rsn20_35 sn20_35 sn21_35 11.551961
Rsp20_36 sp20_36 sp21_36 11.551961
Rsn20_36 sn20_36 sn21_36 11.551961
Rsp20_37 sp20_37 sp21_37 11.551961
Rsn20_37 sn20_37 sn21_37 11.551961
Rsp20_38 sp20_38 sp21_38 11.551961
Rsn20_38 sn20_38 sn21_38 11.551961
Rsp20_39 sp20_39 sp21_39 11.551961
Rsn20_39 sn20_39 sn21_39 11.551961
Rsp20_40 sp20_40 sp21_40 11.551961
Rsn20_40 sn20_40 sn21_40 11.551961
Rsp20_41 sp20_41 sp21_41 11.551961
Rsn20_41 sn20_41 sn21_41 11.551961
Rsp20_42 sp20_42 sp21_42 11.551961
Rsn20_42 sn20_42 sn21_42 11.551961
Rsp20_43 sp20_43 sp21_43 11.551961
Rsn20_43 sn20_43 sn21_43 11.551961
Rsp20_44 sp20_44 sp21_44 11.551961
Rsn20_44 sn20_44 sn21_44 11.551961
Rsp20_45 sp20_45 sp21_45 11.551961
Rsn20_45 sn20_45 sn21_45 11.551961
Rsp20_46 sp20_46 sp21_46 11.551961
Rsn20_46 sn20_46 sn21_46 11.551961
Rsp20_47 sp20_47 sp21_47 11.551961
Rsn20_47 sn20_47 sn21_47 11.551961
Rsp20_48 sp20_48 sp21_48 11.551961
Rsn20_48 sn20_48 sn21_48 11.551961
Rsp20_49 sp20_49 sp21_49 11.551961
Rsn20_49 sn20_49 sn21_49 11.551961
Rsp20_50 sp20_50 sp21_50 11.551961
Rsn20_50 sn20_50 sn21_50 11.551961
Rsp20_51 sp20_51 sp21_51 11.551961
Rsn20_51 sn20_51 sn21_51 11.551961
Rsp20_52 sp20_52 sp21_52 11.551961
Rsn20_52 sn20_52 sn21_52 11.551961
Rsp20_53 sp20_53 sp21_53 11.551961
Rsn20_53 sn20_53 sn21_53 11.551961
Rsp20_54 sp20_54 sp21_54 11.551961
Rsn20_54 sn20_54 sn21_54 11.551961
Rsp20_55 sp20_55 sp21_55 11.551961
Rsn20_55 sn20_55 sn21_55 11.551961
Rsp20_56 sp20_56 sp21_56 11.551961
Rsn20_56 sn20_56 sn21_56 11.551961
Rsp20_57 sp20_57 sp21_57 11.551961
Rsn20_57 sn20_57 sn21_57 11.551961
Rsp20_58 sp20_58 sp21_58 11.551961
Rsn20_58 sn20_58 sn21_58 11.551961
Rsp20_59 sp20_59 sp21_59 11.551961
Rsn20_59 sn20_59 sn21_59 11.551961
Rsp20_60 sp20_60 sp21_60 11.551961
Rsn20_60 sn20_60 sn21_60 11.551961
Rsp20_61 sp20_61 sp21_61 11.551961
Rsn20_61 sn20_61 sn21_61 11.551961
Rsp20_62 sp20_62 sp21_62 11.551961
Rsn20_62 sn20_62 sn21_62 11.551961
Rsp20_63 sp20_63 sp21_63 11.551961
Rsn20_63 sn20_63 sn21_63 11.551961
Rsp20_64 sp20_64 sp21_64 11.551961
Rsn20_64 sn20_64 sn21_64 11.551961
Rsp20_65 sp20_65 sp21_65 11.551961
Rsn20_65 sn20_65 sn21_65 11.551961
Rsp20_66 sp20_66 sp21_66 11.551961
Rsn20_66 sn20_66 sn21_66 11.551961
Rsp20_67 sp20_67 sp21_67 11.551961
Rsn20_67 sn20_67 sn21_67 11.551961
Rsp20_68 sp20_68 sp21_68 11.551961
Rsn20_68 sn20_68 sn21_68 11.551961
Rsp20_69 sp20_69 sp21_69 11.551961
Rsn20_69 sn20_69 sn21_69 11.551961
Rsp20_70 sp20_70 sp21_70 11.551961
Rsn20_70 sn20_70 sn21_70 11.551961
Rsp20_71 sp20_71 sp21_71 11.551961
Rsn20_71 sn20_71 sn21_71 11.551961
Rsp20_72 sp20_72 sp21_72 11.551961
Rsn20_72 sn20_72 sn21_72 11.551961
Rsp20_73 sp20_73 sp21_73 11.551961
Rsn20_73 sn20_73 sn21_73 11.551961
Rsp20_74 sp20_74 sp21_74 11.551961
Rsn20_74 sn20_74 sn21_74 11.551961
Rsp20_75 sp20_75 sp21_75 11.551961
Rsn20_75 sn20_75 sn21_75 11.551961
Rsp20_76 sp20_76 sp21_76 11.551961
Rsn20_76 sn20_76 sn21_76 11.551961
Rsp20_77 sp20_77 sp21_77 11.551961
Rsn20_77 sn20_77 sn21_77 11.551961
Rsp20_78 sp20_78 sp21_78 11.551961
Rsn20_78 sn20_78 sn21_78 11.551961
Rsp20_79 sp20_79 sp21_79 11.551961
Rsn20_79 sn20_79 sn21_79 11.551961
Rsp20_80 sp20_80 sp21_80 11.551961
Rsn20_80 sn20_80 sn21_80 11.551961
Rsp20_81 sp20_81 sp21_81 11.551961
Rsn20_81 sn20_81 sn21_81 11.551961
Rsp20_82 sp20_82 sp21_82 11.551961
Rsn20_82 sn20_82 sn21_82 11.551961
Rsp20_83 sp20_83 sp21_83 11.551961
Rsn20_83 sn20_83 sn21_83 11.551961
Rsp20_84 sp20_84 sp21_84 11.551961
Rsn20_84 sn20_84 sn21_84 11.551961
Rsp21_1 sp21_1 sp22_1 11.551961
Rsn21_1 sn21_1 sn22_1 11.551961
Rsp21_2 sp21_2 sp22_2 11.551961
Rsn21_2 sn21_2 sn22_2 11.551961
Rsp21_3 sp21_3 sp22_3 11.551961
Rsn21_3 sn21_3 sn22_3 11.551961
Rsp21_4 sp21_4 sp22_4 11.551961
Rsn21_4 sn21_4 sn22_4 11.551961
Rsp21_5 sp21_5 sp22_5 11.551961
Rsn21_5 sn21_5 sn22_5 11.551961
Rsp21_6 sp21_6 sp22_6 11.551961
Rsn21_6 sn21_6 sn22_6 11.551961
Rsp21_7 sp21_7 sp22_7 11.551961
Rsn21_7 sn21_7 sn22_7 11.551961
Rsp21_8 sp21_8 sp22_8 11.551961
Rsn21_8 sn21_8 sn22_8 11.551961
Rsp21_9 sp21_9 sp22_9 11.551961
Rsn21_9 sn21_9 sn22_9 11.551961
Rsp21_10 sp21_10 sp22_10 11.551961
Rsn21_10 sn21_10 sn22_10 11.551961
Rsp21_11 sp21_11 sp22_11 11.551961
Rsn21_11 sn21_11 sn22_11 11.551961
Rsp21_12 sp21_12 sp22_12 11.551961
Rsn21_12 sn21_12 sn22_12 11.551961
Rsp21_13 sp21_13 sp22_13 11.551961
Rsn21_13 sn21_13 sn22_13 11.551961
Rsp21_14 sp21_14 sp22_14 11.551961
Rsn21_14 sn21_14 sn22_14 11.551961
Rsp21_15 sp21_15 sp22_15 11.551961
Rsn21_15 sn21_15 sn22_15 11.551961
Rsp21_16 sp21_16 sp22_16 11.551961
Rsn21_16 sn21_16 sn22_16 11.551961
Rsp21_17 sp21_17 sp22_17 11.551961
Rsn21_17 sn21_17 sn22_17 11.551961
Rsp21_18 sp21_18 sp22_18 11.551961
Rsn21_18 sn21_18 sn22_18 11.551961
Rsp21_19 sp21_19 sp22_19 11.551961
Rsn21_19 sn21_19 sn22_19 11.551961
Rsp21_20 sp21_20 sp22_20 11.551961
Rsn21_20 sn21_20 sn22_20 11.551961
Rsp21_21 sp21_21 sp22_21 11.551961
Rsn21_21 sn21_21 sn22_21 11.551961
Rsp21_22 sp21_22 sp22_22 11.551961
Rsn21_22 sn21_22 sn22_22 11.551961
Rsp21_23 sp21_23 sp22_23 11.551961
Rsn21_23 sn21_23 sn22_23 11.551961
Rsp21_24 sp21_24 sp22_24 11.551961
Rsn21_24 sn21_24 sn22_24 11.551961
Rsp21_25 sp21_25 sp22_25 11.551961
Rsn21_25 sn21_25 sn22_25 11.551961
Rsp21_26 sp21_26 sp22_26 11.551961
Rsn21_26 sn21_26 sn22_26 11.551961
Rsp21_27 sp21_27 sp22_27 11.551961
Rsn21_27 sn21_27 sn22_27 11.551961
Rsp21_28 sp21_28 sp22_28 11.551961
Rsn21_28 sn21_28 sn22_28 11.551961
Rsp21_29 sp21_29 sp22_29 11.551961
Rsn21_29 sn21_29 sn22_29 11.551961
Rsp21_30 sp21_30 sp22_30 11.551961
Rsn21_30 sn21_30 sn22_30 11.551961
Rsp21_31 sp21_31 sp22_31 11.551961
Rsn21_31 sn21_31 sn22_31 11.551961
Rsp21_32 sp21_32 sp22_32 11.551961
Rsn21_32 sn21_32 sn22_32 11.551961
Rsp21_33 sp21_33 sp22_33 11.551961
Rsn21_33 sn21_33 sn22_33 11.551961
Rsp21_34 sp21_34 sp22_34 11.551961
Rsn21_34 sn21_34 sn22_34 11.551961
Rsp21_35 sp21_35 sp22_35 11.551961
Rsn21_35 sn21_35 sn22_35 11.551961
Rsp21_36 sp21_36 sp22_36 11.551961
Rsn21_36 sn21_36 sn22_36 11.551961
Rsp21_37 sp21_37 sp22_37 11.551961
Rsn21_37 sn21_37 sn22_37 11.551961
Rsp21_38 sp21_38 sp22_38 11.551961
Rsn21_38 sn21_38 sn22_38 11.551961
Rsp21_39 sp21_39 sp22_39 11.551961
Rsn21_39 sn21_39 sn22_39 11.551961
Rsp21_40 sp21_40 sp22_40 11.551961
Rsn21_40 sn21_40 sn22_40 11.551961
Rsp21_41 sp21_41 sp22_41 11.551961
Rsn21_41 sn21_41 sn22_41 11.551961
Rsp21_42 sp21_42 sp22_42 11.551961
Rsn21_42 sn21_42 sn22_42 11.551961
Rsp21_43 sp21_43 sp22_43 11.551961
Rsn21_43 sn21_43 sn22_43 11.551961
Rsp21_44 sp21_44 sp22_44 11.551961
Rsn21_44 sn21_44 sn22_44 11.551961
Rsp21_45 sp21_45 sp22_45 11.551961
Rsn21_45 sn21_45 sn22_45 11.551961
Rsp21_46 sp21_46 sp22_46 11.551961
Rsn21_46 sn21_46 sn22_46 11.551961
Rsp21_47 sp21_47 sp22_47 11.551961
Rsn21_47 sn21_47 sn22_47 11.551961
Rsp21_48 sp21_48 sp22_48 11.551961
Rsn21_48 sn21_48 sn22_48 11.551961
Rsp21_49 sp21_49 sp22_49 11.551961
Rsn21_49 sn21_49 sn22_49 11.551961
Rsp21_50 sp21_50 sp22_50 11.551961
Rsn21_50 sn21_50 sn22_50 11.551961
Rsp21_51 sp21_51 sp22_51 11.551961
Rsn21_51 sn21_51 sn22_51 11.551961
Rsp21_52 sp21_52 sp22_52 11.551961
Rsn21_52 sn21_52 sn22_52 11.551961
Rsp21_53 sp21_53 sp22_53 11.551961
Rsn21_53 sn21_53 sn22_53 11.551961
Rsp21_54 sp21_54 sp22_54 11.551961
Rsn21_54 sn21_54 sn22_54 11.551961
Rsp21_55 sp21_55 sp22_55 11.551961
Rsn21_55 sn21_55 sn22_55 11.551961
Rsp21_56 sp21_56 sp22_56 11.551961
Rsn21_56 sn21_56 sn22_56 11.551961
Rsp21_57 sp21_57 sp22_57 11.551961
Rsn21_57 sn21_57 sn22_57 11.551961
Rsp21_58 sp21_58 sp22_58 11.551961
Rsn21_58 sn21_58 sn22_58 11.551961
Rsp21_59 sp21_59 sp22_59 11.551961
Rsn21_59 sn21_59 sn22_59 11.551961
Rsp21_60 sp21_60 sp22_60 11.551961
Rsn21_60 sn21_60 sn22_60 11.551961
Rsp21_61 sp21_61 sp22_61 11.551961
Rsn21_61 sn21_61 sn22_61 11.551961
Rsp21_62 sp21_62 sp22_62 11.551961
Rsn21_62 sn21_62 sn22_62 11.551961
Rsp21_63 sp21_63 sp22_63 11.551961
Rsn21_63 sn21_63 sn22_63 11.551961
Rsp21_64 sp21_64 sp22_64 11.551961
Rsn21_64 sn21_64 sn22_64 11.551961
Rsp21_65 sp21_65 sp22_65 11.551961
Rsn21_65 sn21_65 sn22_65 11.551961
Rsp21_66 sp21_66 sp22_66 11.551961
Rsn21_66 sn21_66 sn22_66 11.551961
Rsp21_67 sp21_67 sp22_67 11.551961
Rsn21_67 sn21_67 sn22_67 11.551961
Rsp21_68 sp21_68 sp22_68 11.551961
Rsn21_68 sn21_68 sn22_68 11.551961
Rsp21_69 sp21_69 sp22_69 11.551961
Rsn21_69 sn21_69 sn22_69 11.551961
Rsp21_70 sp21_70 sp22_70 11.551961
Rsn21_70 sn21_70 sn22_70 11.551961
Rsp21_71 sp21_71 sp22_71 11.551961
Rsn21_71 sn21_71 sn22_71 11.551961
Rsp21_72 sp21_72 sp22_72 11.551961
Rsn21_72 sn21_72 sn22_72 11.551961
Rsp21_73 sp21_73 sp22_73 11.551961
Rsn21_73 sn21_73 sn22_73 11.551961
Rsp21_74 sp21_74 sp22_74 11.551961
Rsn21_74 sn21_74 sn22_74 11.551961
Rsp21_75 sp21_75 sp22_75 11.551961
Rsn21_75 sn21_75 sn22_75 11.551961
Rsp21_76 sp21_76 sp22_76 11.551961
Rsn21_76 sn21_76 sn22_76 11.551961
Rsp21_77 sp21_77 sp22_77 11.551961
Rsn21_77 sn21_77 sn22_77 11.551961
Rsp21_78 sp21_78 sp22_78 11.551961
Rsn21_78 sn21_78 sn22_78 11.551961
Rsp21_79 sp21_79 sp22_79 11.551961
Rsn21_79 sn21_79 sn22_79 11.551961
Rsp21_80 sp21_80 sp22_80 11.551961
Rsn21_80 sn21_80 sn22_80 11.551961
Rsp21_81 sp21_81 sp22_81 11.551961
Rsn21_81 sn21_81 sn22_81 11.551961
Rsp21_82 sp21_82 sp22_82 11.551961
Rsn21_82 sn21_82 sn22_82 11.551961
Rsp21_83 sp21_83 sp22_83 11.551961
Rsn21_83 sn21_83 sn22_83 11.551961
Rsp21_84 sp21_84 sp22_84 11.551961
Rsn21_84 sn21_84 sn22_84 11.551961
Rsp22_1 sp22_1 sp23_1 11.551961
Rsn22_1 sn22_1 sn23_1 11.551961
Rsp22_2 sp22_2 sp23_2 11.551961
Rsn22_2 sn22_2 sn23_2 11.551961
Rsp22_3 sp22_3 sp23_3 11.551961
Rsn22_3 sn22_3 sn23_3 11.551961
Rsp22_4 sp22_4 sp23_4 11.551961
Rsn22_4 sn22_4 sn23_4 11.551961
Rsp22_5 sp22_5 sp23_5 11.551961
Rsn22_5 sn22_5 sn23_5 11.551961
Rsp22_6 sp22_6 sp23_6 11.551961
Rsn22_6 sn22_6 sn23_6 11.551961
Rsp22_7 sp22_7 sp23_7 11.551961
Rsn22_7 sn22_7 sn23_7 11.551961
Rsp22_8 sp22_8 sp23_8 11.551961
Rsn22_8 sn22_8 sn23_8 11.551961
Rsp22_9 sp22_9 sp23_9 11.551961
Rsn22_9 sn22_9 sn23_9 11.551961
Rsp22_10 sp22_10 sp23_10 11.551961
Rsn22_10 sn22_10 sn23_10 11.551961
Rsp22_11 sp22_11 sp23_11 11.551961
Rsn22_11 sn22_11 sn23_11 11.551961
Rsp22_12 sp22_12 sp23_12 11.551961
Rsn22_12 sn22_12 sn23_12 11.551961
Rsp22_13 sp22_13 sp23_13 11.551961
Rsn22_13 sn22_13 sn23_13 11.551961
Rsp22_14 sp22_14 sp23_14 11.551961
Rsn22_14 sn22_14 sn23_14 11.551961
Rsp22_15 sp22_15 sp23_15 11.551961
Rsn22_15 sn22_15 sn23_15 11.551961
Rsp22_16 sp22_16 sp23_16 11.551961
Rsn22_16 sn22_16 sn23_16 11.551961
Rsp22_17 sp22_17 sp23_17 11.551961
Rsn22_17 sn22_17 sn23_17 11.551961
Rsp22_18 sp22_18 sp23_18 11.551961
Rsn22_18 sn22_18 sn23_18 11.551961
Rsp22_19 sp22_19 sp23_19 11.551961
Rsn22_19 sn22_19 sn23_19 11.551961
Rsp22_20 sp22_20 sp23_20 11.551961
Rsn22_20 sn22_20 sn23_20 11.551961
Rsp22_21 sp22_21 sp23_21 11.551961
Rsn22_21 sn22_21 sn23_21 11.551961
Rsp22_22 sp22_22 sp23_22 11.551961
Rsn22_22 sn22_22 sn23_22 11.551961
Rsp22_23 sp22_23 sp23_23 11.551961
Rsn22_23 sn22_23 sn23_23 11.551961
Rsp22_24 sp22_24 sp23_24 11.551961
Rsn22_24 sn22_24 sn23_24 11.551961
Rsp22_25 sp22_25 sp23_25 11.551961
Rsn22_25 sn22_25 sn23_25 11.551961
Rsp22_26 sp22_26 sp23_26 11.551961
Rsn22_26 sn22_26 sn23_26 11.551961
Rsp22_27 sp22_27 sp23_27 11.551961
Rsn22_27 sn22_27 sn23_27 11.551961
Rsp22_28 sp22_28 sp23_28 11.551961
Rsn22_28 sn22_28 sn23_28 11.551961
Rsp22_29 sp22_29 sp23_29 11.551961
Rsn22_29 sn22_29 sn23_29 11.551961
Rsp22_30 sp22_30 sp23_30 11.551961
Rsn22_30 sn22_30 sn23_30 11.551961
Rsp22_31 sp22_31 sp23_31 11.551961
Rsn22_31 sn22_31 sn23_31 11.551961
Rsp22_32 sp22_32 sp23_32 11.551961
Rsn22_32 sn22_32 sn23_32 11.551961
Rsp22_33 sp22_33 sp23_33 11.551961
Rsn22_33 sn22_33 sn23_33 11.551961
Rsp22_34 sp22_34 sp23_34 11.551961
Rsn22_34 sn22_34 sn23_34 11.551961
Rsp22_35 sp22_35 sp23_35 11.551961
Rsn22_35 sn22_35 sn23_35 11.551961
Rsp22_36 sp22_36 sp23_36 11.551961
Rsn22_36 sn22_36 sn23_36 11.551961
Rsp22_37 sp22_37 sp23_37 11.551961
Rsn22_37 sn22_37 sn23_37 11.551961
Rsp22_38 sp22_38 sp23_38 11.551961
Rsn22_38 sn22_38 sn23_38 11.551961
Rsp22_39 sp22_39 sp23_39 11.551961
Rsn22_39 sn22_39 sn23_39 11.551961
Rsp22_40 sp22_40 sp23_40 11.551961
Rsn22_40 sn22_40 sn23_40 11.551961
Rsp22_41 sp22_41 sp23_41 11.551961
Rsn22_41 sn22_41 sn23_41 11.551961
Rsp22_42 sp22_42 sp23_42 11.551961
Rsn22_42 sn22_42 sn23_42 11.551961
Rsp22_43 sp22_43 sp23_43 11.551961
Rsn22_43 sn22_43 sn23_43 11.551961
Rsp22_44 sp22_44 sp23_44 11.551961
Rsn22_44 sn22_44 sn23_44 11.551961
Rsp22_45 sp22_45 sp23_45 11.551961
Rsn22_45 sn22_45 sn23_45 11.551961
Rsp22_46 sp22_46 sp23_46 11.551961
Rsn22_46 sn22_46 sn23_46 11.551961
Rsp22_47 sp22_47 sp23_47 11.551961
Rsn22_47 sn22_47 sn23_47 11.551961
Rsp22_48 sp22_48 sp23_48 11.551961
Rsn22_48 sn22_48 sn23_48 11.551961
Rsp22_49 sp22_49 sp23_49 11.551961
Rsn22_49 sn22_49 sn23_49 11.551961
Rsp22_50 sp22_50 sp23_50 11.551961
Rsn22_50 sn22_50 sn23_50 11.551961
Rsp22_51 sp22_51 sp23_51 11.551961
Rsn22_51 sn22_51 sn23_51 11.551961
Rsp22_52 sp22_52 sp23_52 11.551961
Rsn22_52 sn22_52 sn23_52 11.551961
Rsp22_53 sp22_53 sp23_53 11.551961
Rsn22_53 sn22_53 sn23_53 11.551961
Rsp22_54 sp22_54 sp23_54 11.551961
Rsn22_54 sn22_54 sn23_54 11.551961
Rsp22_55 sp22_55 sp23_55 11.551961
Rsn22_55 sn22_55 sn23_55 11.551961
Rsp22_56 sp22_56 sp23_56 11.551961
Rsn22_56 sn22_56 sn23_56 11.551961
Rsp22_57 sp22_57 sp23_57 11.551961
Rsn22_57 sn22_57 sn23_57 11.551961
Rsp22_58 sp22_58 sp23_58 11.551961
Rsn22_58 sn22_58 sn23_58 11.551961
Rsp22_59 sp22_59 sp23_59 11.551961
Rsn22_59 sn22_59 sn23_59 11.551961
Rsp22_60 sp22_60 sp23_60 11.551961
Rsn22_60 sn22_60 sn23_60 11.551961
Rsp22_61 sp22_61 sp23_61 11.551961
Rsn22_61 sn22_61 sn23_61 11.551961
Rsp22_62 sp22_62 sp23_62 11.551961
Rsn22_62 sn22_62 sn23_62 11.551961
Rsp22_63 sp22_63 sp23_63 11.551961
Rsn22_63 sn22_63 sn23_63 11.551961
Rsp22_64 sp22_64 sp23_64 11.551961
Rsn22_64 sn22_64 sn23_64 11.551961
Rsp22_65 sp22_65 sp23_65 11.551961
Rsn22_65 sn22_65 sn23_65 11.551961
Rsp22_66 sp22_66 sp23_66 11.551961
Rsn22_66 sn22_66 sn23_66 11.551961
Rsp22_67 sp22_67 sp23_67 11.551961
Rsn22_67 sn22_67 sn23_67 11.551961
Rsp22_68 sp22_68 sp23_68 11.551961
Rsn22_68 sn22_68 sn23_68 11.551961
Rsp22_69 sp22_69 sp23_69 11.551961
Rsn22_69 sn22_69 sn23_69 11.551961
Rsp22_70 sp22_70 sp23_70 11.551961
Rsn22_70 sn22_70 sn23_70 11.551961
Rsp22_71 sp22_71 sp23_71 11.551961
Rsn22_71 sn22_71 sn23_71 11.551961
Rsp22_72 sp22_72 sp23_72 11.551961
Rsn22_72 sn22_72 sn23_72 11.551961
Rsp22_73 sp22_73 sp23_73 11.551961
Rsn22_73 sn22_73 sn23_73 11.551961
Rsp22_74 sp22_74 sp23_74 11.551961
Rsn22_74 sn22_74 sn23_74 11.551961
Rsp22_75 sp22_75 sp23_75 11.551961
Rsn22_75 sn22_75 sn23_75 11.551961
Rsp22_76 sp22_76 sp23_76 11.551961
Rsn22_76 sn22_76 sn23_76 11.551961
Rsp22_77 sp22_77 sp23_77 11.551961
Rsn22_77 sn22_77 sn23_77 11.551961
Rsp22_78 sp22_78 sp23_78 11.551961
Rsn22_78 sn22_78 sn23_78 11.551961
Rsp22_79 sp22_79 sp23_79 11.551961
Rsn22_79 sn22_79 sn23_79 11.551961
Rsp22_80 sp22_80 sp23_80 11.551961
Rsn22_80 sn22_80 sn23_80 11.551961
Rsp22_81 sp22_81 sp23_81 11.551961
Rsn22_81 sn22_81 sn23_81 11.551961
Rsp22_82 sp22_82 sp23_82 11.551961
Rsn22_82 sn22_82 sn23_82 11.551961
Rsp22_83 sp22_83 sp23_83 11.551961
Rsn22_83 sn22_83 sn23_83 11.551961
Rsp22_84 sp22_84 sp23_84 11.551961
Rsn22_84 sn22_84 sn23_84 11.551961
Rsp23_1 sp23_1 sp24_1 11.551961
Rsn23_1 sn23_1 sn24_1 11.551961
Rsp23_2 sp23_2 sp24_2 11.551961
Rsn23_2 sn23_2 sn24_2 11.551961
Rsp23_3 sp23_3 sp24_3 11.551961
Rsn23_3 sn23_3 sn24_3 11.551961
Rsp23_4 sp23_4 sp24_4 11.551961
Rsn23_4 sn23_4 sn24_4 11.551961
Rsp23_5 sp23_5 sp24_5 11.551961
Rsn23_5 sn23_5 sn24_5 11.551961
Rsp23_6 sp23_6 sp24_6 11.551961
Rsn23_6 sn23_6 sn24_6 11.551961
Rsp23_7 sp23_7 sp24_7 11.551961
Rsn23_7 sn23_7 sn24_7 11.551961
Rsp23_8 sp23_8 sp24_8 11.551961
Rsn23_8 sn23_8 sn24_8 11.551961
Rsp23_9 sp23_9 sp24_9 11.551961
Rsn23_9 sn23_9 sn24_9 11.551961
Rsp23_10 sp23_10 sp24_10 11.551961
Rsn23_10 sn23_10 sn24_10 11.551961
Rsp23_11 sp23_11 sp24_11 11.551961
Rsn23_11 sn23_11 sn24_11 11.551961
Rsp23_12 sp23_12 sp24_12 11.551961
Rsn23_12 sn23_12 sn24_12 11.551961
Rsp23_13 sp23_13 sp24_13 11.551961
Rsn23_13 sn23_13 sn24_13 11.551961
Rsp23_14 sp23_14 sp24_14 11.551961
Rsn23_14 sn23_14 sn24_14 11.551961
Rsp23_15 sp23_15 sp24_15 11.551961
Rsn23_15 sn23_15 sn24_15 11.551961
Rsp23_16 sp23_16 sp24_16 11.551961
Rsn23_16 sn23_16 sn24_16 11.551961
Rsp23_17 sp23_17 sp24_17 11.551961
Rsn23_17 sn23_17 sn24_17 11.551961
Rsp23_18 sp23_18 sp24_18 11.551961
Rsn23_18 sn23_18 sn24_18 11.551961
Rsp23_19 sp23_19 sp24_19 11.551961
Rsn23_19 sn23_19 sn24_19 11.551961
Rsp23_20 sp23_20 sp24_20 11.551961
Rsn23_20 sn23_20 sn24_20 11.551961
Rsp23_21 sp23_21 sp24_21 11.551961
Rsn23_21 sn23_21 sn24_21 11.551961
Rsp23_22 sp23_22 sp24_22 11.551961
Rsn23_22 sn23_22 sn24_22 11.551961
Rsp23_23 sp23_23 sp24_23 11.551961
Rsn23_23 sn23_23 sn24_23 11.551961
Rsp23_24 sp23_24 sp24_24 11.551961
Rsn23_24 sn23_24 sn24_24 11.551961
Rsp23_25 sp23_25 sp24_25 11.551961
Rsn23_25 sn23_25 sn24_25 11.551961
Rsp23_26 sp23_26 sp24_26 11.551961
Rsn23_26 sn23_26 sn24_26 11.551961
Rsp23_27 sp23_27 sp24_27 11.551961
Rsn23_27 sn23_27 sn24_27 11.551961
Rsp23_28 sp23_28 sp24_28 11.551961
Rsn23_28 sn23_28 sn24_28 11.551961
Rsp23_29 sp23_29 sp24_29 11.551961
Rsn23_29 sn23_29 sn24_29 11.551961
Rsp23_30 sp23_30 sp24_30 11.551961
Rsn23_30 sn23_30 sn24_30 11.551961
Rsp23_31 sp23_31 sp24_31 11.551961
Rsn23_31 sn23_31 sn24_31 11.551961
Rsp23_32 sp23_32 sp24_32 11.551961
Rsn23_32 sn23_32 sn24_32 11.551961
Rsp23_33 sp23_33 sp24_33 11.551961
Rsn23_33 sn23_33 sn24_33 11.551961
Rsp23_34 sp23_34 sp24_34 11.551961
Rsn23_34 sn23_34 sn24_34 11.551961
Rsp23_35 sp23_35 sp24_35 11.551961
Rsn23_35 sn23_35 sn24_35 11.551961
Rsp23_36 sp23_36 sp24_36 11.551961
Rsn23_36 sn23_36 sn24_36 11.551961
Rsp23_37 sp23_37 sp24_37 11.551961
Rsn23_37 sn23_37 sn24_37 11.551961
Rsp23_38 sp23_38 sp24_38 11.551961
Rsn23_38 sn23_38 sn24_38 11.551961
Rsp23_39 sp23_39 sp24_39 11.551961
Rsn23_39 sn23_39 sn24_39 11.551961
Rsp23_40 sp23_40 sp24_40 11.551961
Rsn23_40 sn23_40 sn24_40 11.551961
Rsp23_41 sp23_41 sp24_41 11.551961
Rsn23_41 sn23_41 sn24_41 11.551961
Rsp23_42 sp23_42 sp24_42 11.551961
Rsn23_42 sn23_42 sn24_42 11.551961
Rsp23_43 sp23_43 sp24_43 11.551961
Rsn23_43 sn23_43 sn24_43 11.551961
Rsp23_44 sp23_44 sp24_44 11.551961
Rsn23_44 sn23_44 sn24_44 11.551961
Rsp23_45 sp23_45 sp24_45 11.551961
Rsn23_45 sn23_45 sn24_45 11.551961
Rsp23_46 sp23_46 sp24_46 11.551961
Rsn23_46 sn23_46 sn24_46 11.551961
Rsp23_47 sp23_47 sp24_47 11.551961
Rsn23_47 sn23_47 sn24_47 11.551961
Rsp23_48 sp23_48 sp24_48 11.551961
Rsn23_48 sn23_48 sn24_48 11.551961
Rsp23_49 sp23_49 sp24_49 11.551961
Rsn23_49 sn23_49 sn24_49 11.551961
Rsp23_50 sp23_50 sp24_50 11.551961
Rsn23_50 sn23_50 sn24_50 11.551961
Rsp23_51 sp23_51 sp24_51 11.551961
Rsn23_51 sn23_51 sn24_51 11.551961
Rsp23_52 sp23_52 sp24_52 11.551961
Rsn23_52 sn23_52 sn24_52 11.551961
Rsp23_53 sp23_53 sp24_53 11.551961
Rsn23_53 sn23_53 sn24_53 11.551961
Rsp23_54 sp23_54 sp24_54 11.551961
Rsn23_54 sn23_54 sn24_54 11.551961
Rsp23_55 sp23_55 sp24_55 11.551961
Rsn23_55 sn23_55 sn24_55 11.551961
Rsp23_56 sp23_56 sp24_56 11.551961
Rsn23_56 sn23_56 sn24_56 11.551961
Rsp23_57 sp23_57 sp24_57 11.551961
Rsn23_57 sn23_57 sn24_57 11.551961
Rsp23_58 sp23_58 sp24_58 11.551961
Rsn23_58 sn23_58 sn24_58 11.551961
Rsp23_59 sp23_59 sp24_59 11.551961
Rsn23_59 sn23_59 sn24_59 11.551961
Rsp23_60 sp23_60 sp24_60 11.551961
Rsn23_60 sn23_60 sn24_60 11.551961
Rsp23_61 sp23_61 sp24_61 11.551961
Rsn23_61 sn23_61 sn24_61 11.551961
Rsp23_62 sp23_62 sp24_62 11.551961
Rsn23_62 sn23_62 sn24_62 11.551961
Rsp23_63 sp23_63 sp24_63 11.551961
Rsn23_63 sn23_63 sn24_63 11.551961
Rsp23_64 sp23_64 sp24_64 11.551961
Rsn23_64 sn23_64 sn24_64 11.551961
Rsp23_65 sp23_65 sp24_65 11.551961
Rsn23_65 sn23_65 sn24_65 11.551961
Rsp23_66 sp23_66 sp24_66 11.551961
Rsn23_66 sn23_66 sn24_66 11.551961
Rsp23_67 sp23_67 sp24_67 11.551961
Rsn23_67 sn23_67 sn24_67 11.551961
Rsp23_68 sp23_68 sp24_68 11.551961
Rsn23_68 sn23_68 sn24_68 11.551961
Rsp23_69 sp23_69 sp24_69 11.551961
Rsn23_69 sn23_69 sn24_69 11.551961
Rsp23_70 sp23_70 sp24_70 11.551961
Rsn23_70 sn23_70 sn24_70 11.551961
Rsp23_71 sp23_71 sp24_71 11.551961
Rsn23_71 sn23_71 sn24_71 11.551961
Rsp23_72 sp23_72 sp24_72 11.551961
Rsn23_72 sn23_72 sn24_72 11.551961
Rsp23_73 sp23_73 sp24_73 11.551961
Rsn23_73 sn23_73 sn24_73 11.551961
Rsp23_74 sp23_74 sp24_74 11.551961
Rsn23_74 sn23_74 sn24_74 11.551961
Rsp23_75 sp23_75 sp24_75 11.551961
Rsn23_75 sn23_75 sn24_75 11.551961
Rsp23_76 sp23_76 sp24_76 11.551961
Rsn23_76 sn23_76 sn24_76 11.551961
Rsp23_77 sp23_77 sp24_77 11.551961
Rsn23_77 sn23_77 sn24_77 11.551961
Rsp23_78 sp23_78 sp24_78 11.551961
Rsn23_78 sn23_78 sn24_78 11.551961
Rsp23_79 sp23_79 sp24_79 11.551961
Rsn23_79 sn23_79 sn24_79 11.551961
Rsp23_80 sp23_80 sp24_80 11.551961
Rsn23_80 sn23_80 sn24_80 11.551961
Rsp23_81 sp23_81 sp24_81 11.551961
Rsn23_81 sn23_81 sn24_81 11.551961
Rsp23_82 sp23_82 sp24_82 11.551961
Rsn23_82 sn23_82 sn24_82 11.551961
Rsp23_83 sp23_83 sp24_83 11.551961
Rsn23_83 sn23_83 sn24_83 11.551961
Rsp23_84 sp23_84 sp24_84 11.551961
Rsn23_84 sn23_84 sn24_84 11.551961
Rsp24_1 sp24_1 sp25_1 11.551961
Rsn24_1 sn24_1 sn25_1 11.551961
Rsp24_2 sp24_2 sp25_2 11.551961
Rsn24_2 sn24_2 sn25_2 11.551961
Rsp24_3 sp24_3 sp25_3 11.551961
Rsn24_3 sn24_3 sn25_3 11.551961
Rsp24_4 sp24_4 sp25_4 11.551961
Rsn24_4 sn24_4 sn25_4 11.551961
Rsp24_5 sp24_5 sp25_5 11.551961
Rsn24_5 sn24_5 sn25_5 11.551961
Rsp24_6 sp24_6 sp25_6 11.551961
Rsn24_6 sn24_6 sn25_6 11.551961
Rsp24_7 sp24_7 sp25_7 11.551961
Rsn24_7 sn24_7 sn25_7 11.551961
Rsp24_8 sp24_8 sp25_8 11.551961
Rsn24_8 sn24_8 sn25_8 11.551961
Rsp24_9 sp24_9 sp25_9 11.551961
Rsn24_9 sn24_9 sn25_9 11.551961
Rsp24_10 sp24_10 sp25_10 11.551961
Rsn24_10 sn24_10 sn25_10 11.551961
Rsp24_11 sp24_11 sp25_11 11.551961
Rsn24_11 sn24_11 sn25_11 11.551961
Rsp24_12 sp24_12 sp25_12 11.551961
Rsn24_12 sn24_12 sn25_12 11.551961
Rsp24_13 sp24_13 sp25_13 11.551961
Rsn24_13 sn24_13 sn25_13 11.551961
Rsp24_14 sp24_14 sp25_14 11.551961
Rsn24_14 sn24_14 sn25_14 11.551961
Rsp24_15 sp24_15 sp25_15 11.551961
Rsn24_15 sn24_15 sn25_15 11.551961
Rsp24_16 sp24_16 sp25_16 11.551961
Rsn24_16 sn24_16 sn25_16 11.551961
Rsp24_17 sp24_17 sp25_17 11.551961
Rsn24_17 sn24_17 sn25_17 11.551961
Rsp24_18 sp24_18 sp25_18 11.551961
Rsn24_18 sn24_18 sn25_18 11.551961
Rsp24_19 sp24_19 sp25_19 11.551961
Rsn24_19 sn24_19 sn25_19 11.551961
Rsp24_20 sp24_20 sp25_20 11.551961
Rsn24_20 sn24_20 sn25_20 11.551961
Rsp24_21 sp24_21 sp25_21 11.551961
Rsn24_21 sn24_21 sn25_21 11.551961
Rsp24_22 sp24_22 sp25_22 11.551961
Rsn24_22 sn24_22 sn25_22 11.551961
Rsp24_23 sp24_23 sp25_23 11.551961
Rsn24_23 sn24_23 sn25_23 11.551961
Rsp24_24 sp24_24 sp25_24 11.551961
Rsn24_24 sn24_24 sn25_24 11.551961
Rsp24_25 sp24_25 sp25_25 11.551961
Rsn24_25 sn24_25 sn25_25 11.551961
Rsp24_26 sp24_26 sp25_26 11.551961
Rsn24_26 sn24_26 sn25_26 11.551961
Rsp24_27 sp24_27 sp25_27 11.551961
Rsn24_27 sn24_27 sn25_27 11.551961
Rsp24_28 sp24_28 sp25_28 11.551961
Rsn24_28 sn24_28 sn25_28 11.551961
Rsp24_29 sp24_29 sp25_29 11.551961
Rsn24_29 sn24_29 sn25_29 11.551961
Rsp24_30 sp24_30 sp25_30 11.551961
Rsn24_30 sn24_30 sn25_30 11.551961
Rsp24_31 sp24_31 sp25_31 11.551961
Rsn24_31 sn24_31 sn25_31 11.551961
Rsp24_32 sp24_32 sp25_32 11.551961
Rsn24_32 sn24_32 sn25_32 11.551961
Rsp24_33 sp24_33 sp25_33 11.551961
Rsn24_33 sn24_33 sn25_33 11.551961
Rsp24_34 sp24_34 sp25_34 11.551961
Rsn24_34 sn24_34 sn25_34 11.551961
Rsp24_35 sp24_35 sp25_35 11.551961
Rsn24_35 sn24_35 sn25_35 11.551961
Rsp24_36 sp24_36 sp25_36 11.551961
Rsn24_36 sn24_36 sn25_36 11.551961
Rsp24_37 sp24_37 sp25_37 11.551961
Rsn24_37 sn24_37 sn25_37 11.551961
Rsp24_38 sp24_38 sp25_38 11.551961
Rsn24_38 sn24_38 sn25_38 11.551961
Rsp24_39 sp24_39 sp25_39 11.551961
Rsn24_39 sn24_39 sn25_39 11.551961
Rsp24_40 sp24_40 sp25_40 11.551961
Rsn24_40 sn24_40 sn25_40 11.551961
Rsp24_41 sp24_41 sp25_41 11.551961
Rsn24_41 sn24_41 sn25_41 11.551961
Rsp24_42 sp24_42 sp25_42 11.551961
Rsn24_42 sn24_42 sn25_42 11.551961
Rsp24_43 sp24_43 sp25_43 11.551961
Rsn24_43 sn24_43 sn25_43 11.551961
Rsp24_44 sp24_44 sp25_44 11.551961
Rsn24_44 sn24_44 sn25_44 11.551961
Rsp24_45 sp24_45 sp25_45 11.551961
Rsn24_45 sn24_45 sn25_45 11.551961
Rsp24_46 sp24_46 sp25_46 11.551961
Rsn24_46 sn24_46 sn25_46 11.551961
Rsp24_47 sp24_47 sp25_47 11.551961
Rsn24_47 sn24_47 sn25_47 11.551961
Rsp24_48 sp24_48 sp25_48 11.551961
Rsn24_48 sn24_48 sn25_48 11.551961
Rsp24_49 sp24_49 sp25_49 11.551961
Rsn24_49 sn24_49 sn25_49 11.551961
Rsp24_50 sp24_50 sp25_50 11.551961
Rsn24_50 sn24_50 sn25_50 11.551961
Rsp24_51 sp24_51 sp25_51 11.551961
Rsn24_51 sn24_51 sn25_51 11.551961
Rsp24_52 sp24_52 sp25_52 11.551961
Rsn24_52 sn24_52 sn25_52 11.551961
Rsp24_53 sp24_53 sp25_53 11.551961
Rsn24_53 sn24_53 sn25_53 11.551961
Rsp24_54 sp24_54 sp25_54 11.551961
Rsn24_54 sn24_54 sn25_54 11.551961
Rsp24_55 sp24_55 sp25_55 11.551961
Rsn24_55 sn24_55 sn25_55 11.551961
Rsp24_56 sp24_56 sp25_56 11.551961
Rsn24_56 sn24_56 sn25_56 11.551961
Rsp24_57 sp24_57 sp25_57 11.551961
Rsn24_57 sn24_57 sn25_57 11.551961
Rsp24_58 sp24_58 sp25_58 11.551961
Rsn24_58 sn24_58 sn25_58 11.551961
Rsp24_59 sp24_59 sp25_59 11.551961
Rsn24_59 sn24_59 sn25_59 11.551961
Rsp24_60 sp24_60 sp25_60 11.551961
Rsn24_60 sn24_60 sn25_60 11.551961
Rsp24_61 sp24_61 sp25_61 11.551961
Rsn24_61 sn24_61 sn25_61 11.551961
Rsp24_62 sp24_62 sp25_62 11.551961
Rsn24_62 sn24_62 sn25_62 11.551961
Rsp24_63 sp24_63 sp25_63 11.551961
Rsn24_63 sn24_63 sn25_63 11.551961
Rsp24_64 sp24_64 sp25_64 11.551961
Rsn24_64 sn24_64 sn25_64 11.551961
Rsp24_65 sp24_65 sp25_65 11.551961
Rsn24_65 sn24_65 sn25_65 11.551961
Rsp24_66 sp24_66 sp25_66 11.551961
Rsn24_66 sn24_66 sn25_66 11.551961
Rsp24_67 sp24_67 sp25_67 11.551961
Rsn24_67 sn24_67 sn25_67 11.551961
Rsp24_68 sp24_68 sp25_68 11.551961
Rsn24_68 sn24_68 sn25_68 11.551961
Rsp24_69 sp24_69 sp25_69 11.551961
Rsn24_69 sn24_69 sn25_69 11.551961
Rsp24_70 sp24_70 sp25_70 11.551961
Rsn24_70 sn24_70 sn25_70 11.551961
Rsp24_71 sp24_71 sp25_71 11.551961
Rsn24_71 sn24_71 sn25_71 11.551961
Rsp24_72 sp24_72 sp25_72 11.551961
Rsn24_72 sn24_72 sn25_72 11.551961
Rsp24_73 sp24_73 sp25_73 11.551961
Rsn24_73 sn24_73 sn25_73 11.551961
Rsp24_74 sp24_74 sp25_74 11.551961
Rsn24_74 sn24_74 sn25_74 11.551961
Rsp24_75 sp24_75 sp25_75 11.551961
Rsn24_75 sn24_75 sn25_75 11.551961
Rsp24_76 sp24_76 sp25_76 11.551961
Rsn24_76 sn24_76 sn25_76 11.551961
Rsp24_77 sp24_77 sp25_77 11.551961
Rsn24_77 sn24_77 sn25_77 11.551961
Rsp24_78 sp24_78 sp25_78 11.551961
Rsn24_78 sn24_78 sn25_78 11.551961
Rsp24_79 sp24_79 sp25_79 11.551961
Rsn24_79 sn24_79 sn25_79 11.551961
Rsp24_80 sp24_80 sp25_80 11.551961
Rsn24_80 sn24_80 sn25_80 11.551961
Rsp24_81 sp24_81 sp25_81 11.551961
Rsn24_81 sn24_81 sn25_81 11.551961
Rsp24_82 sp24_82 sp25_82 11.551961
Rsn24_82 sn24_82 sn25_82 11.551961
Rsp24_83 sp24_83 sp25_83 11.551961
Rsn24_83 sn24_83 sn25_83 11.551961
Rsp24_84 sp24_84 sp25_84 11.551961
Rsn24_84 sn24_84 sn25_84 11.551961
Rsp25_1 sp25_1 sp26_1 11.551961
Rsn25_1 sn25_1 sn26_1 11.551961
Rsp25_2 sp25_2 sp26_2 11.551961
Rsn25_2 sn25_2 sn26_2 11.551961
Rsp25_3 sp25_3 sp26_3 11.551961
Rsn25_3 sn25_3 sn26_3 11.551961
Rsp25_4 sp25_4 sp26_4 11.551961
Rsn25_4 sn25_4 sn26_4 11.551961
Rsp25_5 sp25_5 sp26_5 11.551961
Rsn25_5 sn25_5 sn26_5 11.551961
Rsp25_6 sp25_6 sp26_6 11.551961
Rsn25_6 sn25_6 sn26_6 11.551961
Rsp25_7 sp25_7 sp26_7 11.551961
Rsn25_7 sn25_7 sn26_7 11.551961
Rsp25_8 sp25_8 sp26_8 11.551961
Rsn25_8 sn25_8 sn26_8 11.551961
Rsp25_9 sp25_9 sp26_9 11.551961
Rsn25_9 sn25_9 sn26_9 11.551961
Rsp25_10 sp25_10 sp26_10 11.551961
Rsn25_10 sn25_10 sn26_10 11.551961
Rsp25_11 sp25_11 sp26_11 11.551961
Rsn25_11 sn25_11 sn26_11 11.551961
Rsp25_12 sp25_12 sp26_12 11.551961
Rsn25_12 sn25_12 sn26_12 11.551961
Rsp25_13 sp25_13 sp26_13 11.551961
Rsn25_13 sn25_13 sn26_13 11.551961
Rsp25_14 sp25_14 sp26_14 11.551961
Rsn25_14 sn25_14 sn26_14 11.551961
Rsp25_15 sp25_15 sp26_15 11.551961
Rsn25_15 sn25_15 sn26_15 11.551961
Rsp25_16 sp25_16 sp26_16 11.551961
Rsn25_16 sn25_16 sn26_16 11.551961
Rsp25_17 sp25_17 sp26_17 11.551961
Rsn25_17 sn25_17 sn26_17 11.551961
Rsp25_18 sp25_18 sp26_18 11.551961
Rsn25_18 sn25_18 sn26_18 11.551961
Rsp25_19 sp25_19 sp26_19 11.551961
Rsn25_19 sn25_19 sn26_19 11.551961
Rsp25_20 sp25_20 sp26_20 11.551961
Rsn25_20 sn25_20 sn26_20 11.551961
Rsp25_21 sp25_21 sp26_21 11.551961
Rsn25_21 sn25_21 sn26_21 11.551961
Rsp25_22 sp25_22 sp26_22 11.551961
Rsn25_22 sn25_22 sn26_22 11.551961
Rsp25_23 sp25_23 sp26_23 11.551961
Rsn25_23 sn25_23 sn26_23 11.551961
Rsp25_24 sp25_24 sp26_24 11.551961
Rsn25_24 sn25_24 sn26_24 11.551961
Rsp25_25 sp25_25 sp26_25 11.551961
Rsn25_25 sn25_25 sn26_25 11.551961
Rsp25_26 sp25_26 sp26_26 11.551961
Rsn25_26 sn25_26 sn26_26 11.551961
Rsp25_27 sp25_27 sp26_27 11.551961
Rsn25_27 sn25_27 sn26_27 11.551961
Rsp25_28 sp25_28 sp26_28 11.551961
Rsn25_28 sn25_28 sn26_28 11.551961
Rsp25_29 sp25_29 sp26_29 11.551961
Rsn25_29 sn25_29 sn26_29 11.551961
Rsp25_30 sp25_30 sp26_30 11.551961
Rsn25_30 sn25_30 sn26_30 11.551961
Rsp25_31 sp25_31 sp26_31 11.551961
Rsn25_31 sn25_31 sn26_31 11.551961
Rsp25_32 sp25_32 sp26_32 11.551961
Rsn25_32 sn25_32 sn26_32 11.551961
Rsp25_33 sp25_33 sp26_33 11.551961
Rsn25_33 sn25_33 sn26_33 11.551961
Rsp25_34 sp25_34 sp26_34 11.551961
Rsn25_34 sn25_34 sn26_34 11.551961
Rsp25_35 sp25_35 sp26_35 11.551961
Rsn25_35 sn25_35 sn26_35 11.551961
Rsp25_36 sp25_36 sp26_36 11.551961
Rsn25_36 sn25_36 sn26_36 11.551961
Rsp25_37 sp25_37 sp26_37 11.551961
Rsn25_37 sn25_37 sn26_37 11.551961
Rsp25_38 sp25_38 sp26_38 11.551961
Rsn25_38 sn25_38 sn26_38 11.551961
Rsp25_39 sp25_39 sp26_39 11.551961
Rsn25_39 sn25_39 sn26_39 11.551961
Rsp25_40 sp25_40 sp26_40 11.551961
Rsn25_40 sn25_40 sn26_40 11.551961
Rsp25_41 sp25_41 sp26_41 11.551961
Rsn25_41 sn25_41 sn26_41 11.551961
Rsp25_42 sp25_42 sp26_42 11.551961
Rsn25_42 sn25_42 sn26_42 11.551961
Rsp25_43 sp25_43 sp26_43 11.551961
Rsn25_43 sn25_43 sn26_43 11.551961
Rsp25_44 sp25_44 sp26_44 11.551961
Rsn25_44 sn25_44 sn26_44 11.551961
Rsp25_45 sp25_45 sp26_45 11.551961
Rsn25_45 sn25_45 sn26_45 11.551961
Rsp25_46 sp25_46 sp26_46 11.551961
Rsn25_46 sn25_46 sn26_46 11.551961
Rsp25_47 sp25_47 sp26_47 11.551961
Rsn25_47 sn25_47 sn26_47 11.551961
Rsp25_48 sp25_48 sp26_48 11.551961
Rsn25_48 sn25_48 sn26_48 11.551961
Rsp25_49 sp25_49 sp26_49 11.551961
Rsn25_49 sn25_49 sn26_49 11.551961
Rsp25_50 sp25_50 sp26_50 11.551961
Rsn25_50 sn25_50 sn26_50 11.551961
Rsp25_51 sp25_51 sp26_51 11.551961
Rsn25_51 sn25_51 sn26_51 11.551961
Rsp25_52 sp25_52 sp26_52 11.551961
Rsn25_52 sn25_52 sn26_52 11.551961
Rsp25_53 sp25_53 sp26_53 11.551961
Rsn25_53 sn25_53 sn26_53 11.551961
Rsp25_54 sp25_54 sp26_54 11.551961
Rsn25_54 sn25_54 sn26_54 11.551961
Rsp25_55 sp25_55 sp26_55 11.551961
Rsn25_55 sn25_55 sn26_55 11.551961
Rsp25_56 sp25_56 sp26_56 11.551961
Rsn25_56 sn25_56 sn26_56 11.551961
Rsp25_57 sp25_57 sp26_57 11.551961
Rsn25_57 sn25_57 sn26_57 11.551961
Rsp25_58 sp25_58 sp26_58 11.551961
Rsn25_58 sn25_58 sn26_58 11.551961
Rsp25_59 sp25_59 sp26_59 11.551961
Rsn25_59 sn25_59 sn26_59 11.551961
Rsp25_60 sp25_60 sp26_60 11.551961
Rsn25_60 sn25_60 sn26_60 11.551961
Rsp25_61 sp25_61 sp26_61 11.551961
Rsn25_61 sn25_61 sn26_61 11.551961
Rsp25_62 sp25_62 sp26_62 11.551961
Rsn25_62 sn25_62 sn26_62 11.551961
Rsp25_63 sp25_63 sp26_63 11.551961
Rsn25_63 sn25_63 sn26_63 11.551961
Rsp25_64 sp25_64 sp26_64 11.551961
Rsn25_64 sn25_64 sn26_64 11.551961
Rsp25_65 sp25_65 sp26_65 11.551961
Rsn25_65 sn25_65 sn26_65 11.551961
Rsp25_66 sp25_66 sp26_66 11.551961
Rsn25_66 sn25_66 sn26_66 11.551961
Rsp25_67 sp25_67 sp26_67 11.551961
Rsn25_67 sn25_67 sn26_67 11.551961
Rsp25_68 sp25_68 sp26_68 11.551961
Rsn25_68 sn25_68 sn26_68 11.551961
Rsp25_69 sp25_69 sp26_69 11.551961
Rsn25_69 sn25_69 sn26_69 11.551961
Rsp25_70 sp25_70 sp26_70 11.551961
Rsn25_70 sn25_70 sn26_70 11.551961
Rsp25_71 sp25_71 sp26_71 11.551961
Rsn25_71 sn25_71 sn26_71 11.551961
Rsp25_72 sp25_72 sp26_72 11.551961
Rsn25_72 sn25_72 sn26_72 11.551961
Rsp25_73 sp25_73 sp26_73 11.551961
Rsn25_73 sn25_73 sn26_73 11.551961
Rsp25_74 sp25_74 sp26_74 11.551961
Rsn25_74 sn25_74 sn26_74 11.551961
Rsp25_75 sp25_75 sp26_75 11.551961
Rsn25_75 sn25_75 sn26_75 11.551961
Rsp25_76 sp25_76 sp26_76 11.551961
Rsn25_76 sn25_76 sn26_76 11.551961
Rsp25_77 sp25_77 sp26_77 11.551961
Rsn25_77 sn25_77 sn26_77 11.551961
Rsp25_78 sp25_78 sp26_78 11.551961
Rsn25_78 sn25_78 sn26_78 11.551961
Rsp25_79 sp25_79 sp26_79 11.551961
Rsn25_79 sn25_79 sn26_79 11.551961
Rsp25_80 sp25_80 sp26_80 11.551961
Rsn25_80 sn25_80 sn26_80 11.551961
Rsp25_81 sp25_81 sp26_81 11.551961
Rsn25_81 sn25_81 sn26_81 11.551961
Rsp25_82 sp25_82 sp26_82 11.551961
Rsn25_82 sn25_82 sn26_82 11.551961
Rsp25_83 sp25_83 sp26_83 11.551961
Rsn25_83 sn25_83 sn26_83 11.551961
Rsp25_84 sp25_84 sp26_84 11.551961
Rsn25_84 sn25_84 sn26_84 11.551961
Rsp26_1 sp26_1 sp27_1 11.551961
Rsn26_1 sn26_1 sn27_1 11.551961
Rsp26_2 sp26_2 sp27_2 11.551961
Rsn26_2 sn26_2 sn27_2 11.551961
Rsp26_3 sp26_3 sp27_3 11.551961
Rsn26_3 sn26_3 sn27_3 11.551961
Rsp26_4 sp26_4 sp27_4 11.551961
Rsn26_4 sn26_4 sn27_4 11.551961
Rsp26_5 sp26_5 sp27_5 11.551961
Rsn26_5 sn26_5 sn27_5 11.551961
Rsp26_6 sp26_6 sp27_6 11.551961
Rsn26_6 sn26_6 sn27_6 11.551961
Rsp26_7 sp26_7 sp27_7 11.551961
Rsn26_7 sn26_7 sn27_7 11.551961
Rsp26_8 sp26_8 sp27_8 11.551961
Rsn26_8 sn26_8 sn27_8 11.551961
Rsp26_9 sp26_9 sp27_9 11.551961
Rsn26_9 sn26_9 sn27_9 11.551961
Rsp26_10 sp26_10 sp27_10 11.551961
Rsn26_10 sn26_10 sn27_10 11.551961
Rsp26_11 sp26_11 sp27_11 11.551961
Rsn26_11 sn26_11 sn27_11 11.551961
Rsp26_12 sp26_12 sp27_12 11.551961
Rsn26_12 sn26_12 sn27_12 11.551961
Rsp26_13 sp26_13 sp27_13 11.551961
Rsn26_13 sn26_13 sn27_13 11.551961
Rsp26_14 sp26_14 sp27_14 11.551961
Rsn26_14 sn26_14 sn27_14 11.551961
Rsp26_15 sp26_15 sp27_15 11.551961
Rsn26_15 sn26_15 sn27_15 11.551961
Rsp26_16 sp26_16 sp27_16 11.551961
Rsn26_16 sn26_16 sn27_16 11.551961
Rsp26_17 sp26_17 sp27_17 11.551961
Rsn26_17 sn26_17 sn27_17 11.551961
Rsp26_18 sp26_18 sp27_18 11.551961
Rsn26_18 sn26_18 sn27_18 11.551961
Rsp26_19 sp26_19 sp27_19 11.551961
Rsn26_19 sn26_19 sn27_19 11.551961
Rsp26_20 sp26_20 sp27_20 11.551961
Rsn26_20 sn26_20 sn27_20 11.551961
Rsp26_21 sp26_21 sp27_21 11.551961
Rsn26_21 sn26_21 sn27_21 11.551961
Rsp26_22 sp26_22 sp27_22 11.551961
Rsn26_22 sn26_22 sn27_22 11.551961
Rsp26_23 sp26_23 sp27_23 11.551961
Rsn26_23 sn26_23 sn27_23 11.551961
Rsp26_24 sp26_24 sp27_24 11.551961
Rsn26_24 sn26_24 sn27_24 11.551961
Rsp26_25 sp26_25 sp27_25 11.551961
Rsn26_25 sn26_25 sn27_25 11.551961
Rsp26_26 sp26_26 sp27_26 11.551961
Rsn26_26 sn26_26 sn27_26 11.551961
Rsp26_27 sp26_27 sp27_27 11.551961
Rsn26_27 sn26_27 sn27_27 11.551961
Rsp26_28 sp26_28 sp27_28 11.551961
Rsn26_28 sn26_28 sn27_28 11.551961
Rsp26_29 sp26_29 sp27_29 11.551961
Rsn26_29 sn26_29 sn27_29 11.551961
Rsp26_30 sp26_30 sp27_30 11.551961
Rsn26_30 sn26_30 sn27_30 11.551961
Rsp26_31 sp26_31 sp27_31 11.551961
Rsn26_31 sn26_31 sn27_31 11.551961
Rsp26_32 sp26_32 sp27_32 11.551961
Rsn26_32 sn26_32 sn27_32 11.551961
Rsp26_33 sp26_33 sp27_33 11.551961
Rsn26_33 sn26_33 sn27_33 11.551961
Rsp26_34 sp26_34 sp27_34 11.551961
Rsn26_34 sn26_34 sn27_34 11.551961
Rsp26_35 sp26_35 sp27_35 11.551961
Rsn26_35 sn26_35 sn27_35 11.551961
Rsp26_36 sp26_36 sp27_36 11.551961
Rsn26_36 sn26_36 sn27_36 11.551961
Rsp26_37 sp26_37 sp27_37 11.551961
Rsn26_37 sn26_37 sn27_37 11.551961
Rsp26_38 sp26_38 sp27_38 11.551961
Rsn26_38 sn26_38 sn27_38 11.551961
Rsp26_39 sp26_39 sp27_39 11.551961
Rsn26_39 sn26_39 sn27_39 11.551961
Rsp26_40 sp26_40 sp27_40 11.551961
Rsn26_40 sn26_40 sn27_40 11.551961
Rsp26_41 sp26_41 sp27_41 11.551961
Rsn26_41 sn26_41 sn27_41 11.551961
Rsp26_42 sp26_42 sp27_42 11.551961
Rsn26_42 sn26_42 sn27_42 11.551961
Rsp26_43 sp26_43 sp27_43 11.551961
Rsn26_43 sn26_43 sn27_43 11.551961
Rsp26_44 sp26_44 sp27_44 11.551961
Rsn26_44 sn26_44 sn27_44 11.551961
Rsp26_45 sp26_45 sp27_45 11.551961
Rsn26_45 sn26_45 sn27_45 11.551961
Rsp26_46 sp26_46 sp27_46 11.551961
Rsn26_46 sn26_46 sn27_46 11.551961
Rsp26_47 sp26_47 sp27_47 11.551961
Rsn26_47 sn26_47 sn27_47 11.551961
Rsp26_48 sp26_48 sp27_48 11.551961
Rsn26_48 sn26_48 sn27_48 11.551961
Rsp26_49 sp26_49 sp27_49 11.551961
Rsn26_49 sn26_49 sn27_49 11.551961
Rsp26_50 sp26_50 sp27_50 11.551961
Rsn26_50 sn26_50 sn27_50 11.551961
Rsp26_51 sp26_51 sp27_51 11.551961
Rsn26_51 sn26_51 sn27_51 11.551961
Rsp26_52 sp26_52 sp27_52 11.551961
Rsn26_52 sn26_52 sn27_52 11.551961
Rsp26_53 sp26_53 sp27_53 11.551961
Rsn26_53 sn26_53 sn27_53 11.551961
Rsp26_54 sp26_54 sp27_54 11.551961
Rsn26_54 sn26_54 sn27_54 11.551961
Rsp26_55 sp26_55 sp27_55 11.551961
Rsn26_55 sn26_55 sn27_55 11.551961
Rsp26_56 sp26_56 sp27_56 11.551961
Rsn26_56 sn26_56 sn27_56 11.551961
Rsp26_57 sp26_57 sp27_57 11.551961
Rsn26_57 sn26_57 sn27_57 11.551961
Rsp26_58 sp26_58 sp27_58 11.551961
Rsn26_58 sn26_58 sn27_58 11.551961
Rsp26_59 sp26_59 sp27_59 11.551961
Rsn26_59 sn26_59 sn27_59 11.551961
Rsp26_60 sp26_60 sp27_60 11.551961
Rsn26_60 sn26_60 sn27_60 11.551961
Rsp26_61 sp26_61 sp27_61 11.551961
Rsn26_61 sn26_61 sn27_61 11.551961
Rsp26_62 sp26_62 sp27_62 11.551961
Rsn26_62 sn26_62 sn27_62 11.551961
Rsp26_63 sp26_63 sp27_63 11.551961
Rsn26_63 sn26_63 sn27_63 11.551961
Rsp26_64 sp26_64 sp27_64 11.551961
Rsn26_64 sn26_64 sn27_64 11.551961
Rsp26_65 sp26_65 sp27_65 11.551961
Rsn26_65 sn26_65 sn27_65 11.551961
Rsp26_66 sp26_66 sp27_66 11.551961
Rsn26_66 sn26_66 sn27_66 11.551961
Rsp26_67 sp26_67 sp27_67 11.551961
Rsn26_67 sn26_67 sn27_67 11.551961
Rsp26_68 sp26_68 sp27_68 11.551961
Rsn26_68 sn26_68 sn27_68 11.551961
Rsp26_69 sp26_69 sp27_69 11.551961
Rsn26_69 sn26_69 sn27_69 11.551961
Rsp26_70 sp26_70 sp27_70 11.551961
Rsn26_70 sn26_70 sn27_70 11.551961
Rsp26_71 sp26_71 sp27_71 11.551961
Rsn26_71 sn26_71 sn27_71 11.551961
Rsp26_72 sp26_72 sp27_72 11.551961
Rsn26_72 sn26_72 sn27_72 11.551961
Rsp26_73 sp26_73 sp27_73 11.551961
Rsn26_73 sn26_73 sn27_73 11.551961
Rsp26_74 sp26_74 sp27_74 11.551961
Rsn26_74 sn26_74 sn27_74 11.551961
Rsp26_75 sp26_75 sp27_75 11.551961
Rsn26_75 sn26_75 sn27_75 11.551961
Rsp26_76 sp26_76 sp27_76 11.551961
Rsn26_76 sn26_76 sn27_76 11.551961
Rsp26_77 sp26_77 sp27_77 11.551961
Rsn26_77 sn26_77 sn27_77 11.551961
Rsp26_78 sp26_78 sp27_78 11.551961
Rsn26_78 sn26_78 sn27_78 11.551961
Rsp26_79 sp26_79 sp27_79 11.551961
Rsn26_79 sn26_79 sn27_79 11.551961
Rsp26_80 sp26_80 sp27_80 11.551961
Rsn26_80 sn26_80 sn27_80 11.551961
Rsp26_81 sp26_81 sp27_81 11.551961
Rsn26_81 sn26_81 sn27_81 11.551961
Rsp26_82 sp26_82 sp27_82 11.551961
Rsn26_82 sn26_82 sn27_82 11.551961
Rsp26_83 sp26_83 sp27_83 11.551961
Rsn26_83 sn26_83 sn27_83 11.551961
Rsp26_84 sp26_84 sp27_84 11.551961
Rsn26_84 sn26_84 sn27_84 11.551961
Rsp27_1 sp27_1 sp28_1 11.551961
Rsn27_1 sn27_1 sn28_1 11.551961
Rsp27_2 sp27_2 sp28_2 11.551961
Rsn27_2 sn27_2 sn28_2 11.551961
Rsp27_3 sp27_3 sp28_3 11.551961
Rsn27_3 sn27_3 sn28_3 11.551961
Rsp27_4 sp27_4 sp28_4 11.551961
Rsn27_4 sn27_4 sn28_4 11.551961
Rsp27_5 sp27_5 sp28_5 11.551961
Rsn27_5 sn27_5 sn28_5 11.551961
Rsp27_6 sp27_6 sp28_6 11.551961
Rsn27_6 sn27_6 sn28_6 11.551961
Rsp27_7 sp27_7 sp28_7 11.551961
Rsn27_7 sn27_7 sn28_7 11.551961
Rsp27_8 sp27_8 sp28_8 11.551961
Rsn27_8 sn27_8 sn28_8 11.551961
Rsp27_9 sp27_9 sp28_9 11.551961
Rsn27_9 sn27_9 sn28_9 11.551961
Rsp27_10 sp27_10 sp28_10 11.551961
Rsn27_10 sn27_10 sn28_10 11.551961
Rsp27_11 sp27_11 sp28_11 11.551961
Rsn27_11 sn27_11 sn28_11 11.551961
Rsp27_12 sp27_12 sp28_12 11.551961
Rsn27_12 sn27_12 sn28_12 11.551961
Rsp27_13 sp27_13 sp28_13 11.551961
Rsn27_13 sn27_13 sn28_13 11.551961
Rsp27_14 sp27_14 sp28_14 11.551961
Rsn27_14 sn27_14 sn28_14 11.551961
Rsp27_15 sp27_15 sp28_15 11.551961
Rsn27_15 sn27_15 sn28_15 11.551961
Rsp27_16 sp27_16 sp28_16 11.551961
Rsn27_16 sn27_16 sn28_16 11.551961
Rsp27_17 sp27_17 sp28_17 11.551961
Rsn27_17 sn27_17 sn28_17 11.551961
Rsp27_18 sp27_18 sp28_18 11.551961
Rsn27_18 sn27_18 sn28_18 11.551961
Rsp27_19 sp27_19 sp28_19 11.551961
Rsn27_19 sn27_19 sn28_19 11.551961
Rsp27_20 sp27_20 sp28_20 11.551961
Rsn27_20 sn27_20 sn28_20 11.551961
Rsp27_21 sp27_21 sp28_21 11.551961
Rsn27_21 sn27_21 sn28_21 11.551961
Rsp27_22 sp27_22 sp28_22 11.551961
Rsn27_22 sn27_22 sn28_22 11.551961
Rsp27_23 sp27_23 sp28_23 11.551961
Rsn27_23 sn27_23 sn28_23 11.551961
Rsp27_24 sp27_24 sp28_24 11.551961
Rsn27_24 sn27_24 sn28_24 11.551961
Rsp27_25 sp27_25 sp28_25 11.551961
Rsn27_25 sn27_25 sn28_25 11.551961
Rsp27_26 sp27_26 sp28_26 11.551961
Rsn27_26 sn27_26 sn28_26 11.551961
Rsp27_27 sp27_27 sp28_27 11.551961
Rsn27_27 sn27_27 sn28_27 11.551961
Rsp27_28 sp27_28 sp28_28 11.551961
Rsn27_28 sn27_28 sn28_28 11.551961
Rsp27_29 sp27_29 sp28_29 11.551961
Rsn27_29 sn27_29 sn28_29 11.551961
Rsp27_30 sp27_30 sp28_30 11.551961
Rsn27_30 sn27_30 sn28_30 11.551961
Rsp27_31 sp27_31 sp28_31 11.551961
Rsn27_31 sn27_31 sn28_31 11.551961
Rsp27_32 sp27_32 sp28_32 11.551961
Rsn27_32 sn27_32 sn28_32 11.551961
Rsp27_33 sp27_33 sp28_33 11.551961
Rsn27_33 sn27_33 sn28_33 11.551961
Rsp27_34 sp27_34 sp28_34 11.551961
Rsn27_34 sn27_34 sn28_34 11.551961
Rsp27_35 sp27_35 sp28_35 11.551961
Rsn27_35 sn27_35 sn28_35 11.551961
Rsp27_36 sp27_36 sp28_36 11.551961
Rsn27_36 sn27_36 sn28_36 11.551961
Rsp27_37 sp27_37 sp28_37 11.551961
Rsn27_37 sn27_37 sn28_37 11.551961
Rsp27_38 sp27_38 sp28_38 11.551961
Rsn27_38 sn27_38 sn28_38 11.551961
Rsp27_39 sp27_39 sp28_39 11.551961
Rsn27_39 sn27_39 sn28_39 11.551961
Rsp27_40 sp27_40 sp28_40 11.551961
Rsn27_40 sn27_40 sn28_40 11.551961
Rsp27_41 sp27_41 sp28_41 11.551961
Rsn27_41 sn27_41 sn28_41 11.551961
Rsp27_42 sp27_42 sp28_42 11.551961
Rsn27_42 sn27_42 sn28_42 11.551961
Rsp27_43 sp27_43 sp28_43 11.551961
Rsn27_43 sn27_43 sn28_43 11.551961
Rsp27_44 sp27_44 sp28_44 11.551961
Rsn27_44 sn27_44 sn28_44 11.551961
Rsp27_45 sp27_45 sp28_45 11.551961
Rsn27_45 sn27_45 sn28_45 11.551961
Rsp27_46 sp27_46 sp28_46 11.551961
Rsn27_46 sn27_46 sn28_46 11.551961
Rsp27_47 sp27_47 sp28_47 11.551961
Rsn27_47 sn27_47 sn28_47 11.551961
Rsp27_48 sp27_48 sp28_48 11.551961
Rsn27_48 sn27_48 sn28_48 11.551961
Rsp27_49 sp27_49 sp28_49 11.551961
Rsn27_49 sn27_49 sn28_49 11.551961
Rsp27_50 sp27_50 sp28_50 11.551961
Rsn27_50 sn27_50 sn28_50 11.551961
Rsp27_51 sp27_51 sp28_51 11.551961
Rsn27_51 sn27_51 sn28_51 11.551961
Rsp27_52 sp27_52 sp28_52 11.551961
Rsn27_52 sn27_52 sn28_52 11.551961
Rsp27_53 sp27_53 sp28_53 11.551961
Rsn27_53 sn27_53 sn28_53 11.551961
Rsp27_54 sp27_54 sp28_54 11.551961
Rsn27_54 sn27_54 sn28_54 11.551961
Rsp27_55 sp27_55 sp28_55 11.551961
Rsn27_55 sn27_55 sn28_55 11.551961
Rsp27_56 sp27_56 sp28_56 11.551961
Rsn27_56 sn27_56 sn28_56 11.551961
Rsp27_57 sp27_57 sp28_57 11.551961
Rsn27_57 sn27_57 sn28_57 11.551961
Rsp27_58 sp27_58 sp28_58 11.551961
Rsn27_58 sn27_58 sn28_58 11.551961
Rsp27_59 sp27_59 sp28_59 11.551961
Rsn27_59 sn27_59 sn28_59 11.551961
Rsp27_60 sp27_60 sp28_60 11.551961
Rsn27_60 sn27_60 sn28_60 11.551961
Rsp27_61 sp27_61 sp28_61 11.551961
Rsn27_61 sn27_61 sn28_61 11.551961
Rsp27_62 sp27_62 sp28_62 11.551961
Rsn27_62 sn27_62 sn28_62 11.551961
Rsp27_63 sp27_63 sp28_63 11.551961
Rsn27_63 sn27_63 sn28_63 11.551961
Rsp27_64 sp27_64 sp28_64 11.551961
Rsn27_64 sn27_64 sn28_64 11.551961
Rsp27_65 sp27_65 sp28_65 11.551961
Rsn27_65 sn27_65 sn28_65 11.551961
Rsp27_66 sp27_66 sp28_66 11.551961
Rsn27_66 sn27_66 sn28_66 11.551961
Rsp27_67 sp27_67 sp28_67 11.551961
Rsn27_67 sn27_67 sn28_67 11.551961
Rsp27_68 sp27_68 sp28_68 11.551961
Rsn27_68 sn27_68 sn28_68 11.551961
Rsp27_69 sp27_69 sp28_69 11.551961
Rsn27_69 sn27_69 sn28_69 11.551961
Rsp27_70 sp27_70 sp28_70 11.551961
Rsn27_70 sn27_70 sn28_70 11.551961
Rsp27_71 sp27_71 sp28_71 11.551961
Rsn27_71 sn27_71 sn28_71 11.551961
Rsp27_72 sp27_72 sp28_72 11.551961
Rsn27_72 sn27_72 sn28_72 11.551961
Rsp27_73 sp27_73 sp28_73 11.551961
Rsn27_73 sn27_73 sn28_73 11.551961
Rsp27_74 sp27_74 sp28_74 11.551961
Rsn27_74 sn27_74 sn28_74 11.551961
Rsp27_75 sp27_75 sp28_75 11.551961
Rsn27_75 sn27_75 sn28_75 11.551961
Rsp27_76 sp27_76 sp28_76 11.551961
Rsn27_76 sn27_76 sn28_76 11.551961
Rsp27_77 sp27_77 sp28_77 11.551961
Rsn27_77 sn27_77 sn28_77 11.551961
Rsp27_78 sp27_78 sp28_78 11.551961
Rsn27_78 sn27_78 sn28_78 11.551961
Rsp27_79 sp27_79 sp28_79 11.551961
Rsn27_79 sn27_79 sn28_79 11.551961
Rsp27_80 sp27_80 sp28_80 11.551961
Rsn27_80 sn27_80 sn28_80 11.551961
Rsp27_81 sp27_81 sp28_81 11.551961
Rsn27_81 sn27_81 sn28_81 11.551961
Rsp27_82 sp27_82 sp28_82 11.551961
Rsn27_82 sn27_82 sn28_82 11.551961
Rsp27_83 sp27_83 sp28_83 11.551961
Rsn27_83 sn27_83 sn28_83 11.551961
Rsp27_84 sp27_84 sp28_84 11.551961
Rsn27_84 sn27_84 sn28_84 11.551961
Rsp28_1 sp28_1 sp29_1 11.551961
Rsn28_1 sn28_1 sn29_1 11.551961
Rsp28_2 sp28_2 sp29_2 11.551961
Rsn28_2 sn28_2 sn29_2 11.551961
Rsp28_3 sp28_3 sp29_3 11.551961
Rsn28_3 sn28_3 sn29_3 11.551961
Rsp28_4 sp28_4 sp29_4 11.551961
Rsn28_4 sn28_4 sn29_4 11.551961
Rsp28_5 sp28_5 sp29_5 11.551961
Rsn28_5 sn28_5 sn29_5 11.551961
Rsp28_6 sp28_6 sp29_6 11.551961
Rsn28_6 sn28_6 sn29_6 11.551961
Rsp28_7 sp28_7 sp29_7 11.551961
Rsn28_7 sn28_7 sn29_7 11.551961
Rsp28_8 sp28_8 sp29_8 11.551961
Rsn28_8 sn28_8 sn29_8 11.551961
Rsp28_9 sp28_9 sp29_9 11.551961
Rsn28_9 sn28_9 sn29_9 11.551961
Rsp28_10 sp28_10 sp29_10 11.551961
Rsn28_10 sn28_10 sn29_10 11.551961
Rsp28_11 sp28_11 sp29_11 11.551961
Rsn28_11 sn28_11 sn29_11 11.551961
Rsp28_12 sp28_12 sp29_12 11.551961
Rsn28_12 sn28_12 sn29_12 11.551961
Rsp28_13 sp28_13 sp29_13 11.551961
Rsn28_13 sn28_13 sn29_13 11.551961
Rsp28_14 sp28_14 sp29_14 11.551961
Rsn28_14 sn28_14 sn29_14 11.551961
Rsp28_15 sp28_15 sp29_15 11.551961
Rsn28_15 sn28_15 sn29_15 11.551961
Rsp28_16 sp28_16 sp29_16 11.551961
Rsn28_16 sn28_16 sn29_16 11.551961
Rsp28_17 sp28_17 sp29_17 11.551961
Rsn28_17 sn28_17 sn29_17 11.551961
Rsp28_18 sp28_18 sp29_18 11.551961
Rsn28_18 sn28_18 sn29_18 11.551961
Rsp28_19 sp28_19 sp29_19 11.551961
Rsn28_19 sn28_19 sn29_19 11.551961
Rsp28_20 sp28_20 sp29_20 11.551961
Rsn28_20 sn28_20 sn29_20 11.551961
Rsp28_21 sp28_21 sp29_21 11.551961
Rsn28_21 sn28_21 sn29_21 11.551961
Rsp28_22 sp28_22 sp29_22 11.551961
Rsn28_22 sn28_22 sn29_22 11.551961
Rsp28_23 sp28_23 sp29_23 11.551961
Rsn28_23 sn28_23 sn29_23 11.551961
Rsp28_24 sp28_24 sp29_24 11.551961
Rsn28_24 sn28_24 sn29_24 11.551961
Rsp28_25 sp28_25 sp29_25 11.551961
Rsn28_25 sn28_25 sn29_25 11.551961
Rsp28_26 sp28_26 sp29_26 11.551961
Rsn28_26 sn28_26 sn29_26 11.551961
Rsp28_27 sp28_27 sp29_27 11.551961
Rsn28_27 sn28_27 sn29_27 11.551961
Rsp28_28 sp28_28 sp29_28 11.551961
Rsn28_28 sn28_28 sn29_28 11.551961
Rsp28_29 sp28_29 sp29_29 11.551961
Rsn28_29 sn28_29 sn29_29 11.551961
Rsp28_30 sp28_30 sp29_30 11.551961
Rsn28_30 sn28_30 sn29_30 11.551961
Rsp28_31 sp28_31 sp29_31 11.551961
Rsn28_31 sn28_31 sn29_31 11.551961
Rsp28_32 sp28_32 sp29_32 11.551961
Rsn28_32 sn28_32 sn29_32 11.551961
Rsp28_33 sp28_33 sp29_33 11.551961
Rsn28_33 sn28_33 sn29_33 11.551961
Rsp28_34 sp28_34 sp29_34 11.551961
Rsn28_34 sn28_34 sn29_34 11.551961
Rsp28_35 sp28_35 sp29_35 11.551961
Rsn28_35 sn28_35 sn29_35 11.551961
Rsp28_36 sp28_36 sp29_36 11.551961
Rsn28_36 sn28_36 sn29_36 11.551961
Rsp28_37 sp28_37 sp29_37 11.551961
Rsn28_37 sn28_37 sn29_37 11.551961
Rsp28_38 sp28_38 sp29_38 11.551961
Rsn28_38 sn28_38 sn29_38 11.551961
Rsp28_39 sp28_39 sp29_39 11.551961
Rsn28_39 sn28_39 sn29_39 11.551961
Rsp28_40 sp28_40 sp29_40 11.551961
Rsn28_40 sn28_40 sn29_40 11.551961
Rsp28_41 sp28_41 sp29_41 11.551961
Rsn28_41 sn28_41 sn29_41 11.551961
Rsp28_42 sp28_42 sp29_42 11.551961
Rsn28_42 sn28_42 sn29_42 11.551961
Rsp28_43 sp28_43 sp29_43 11.551961
Rsn28_43 sn28_43 sn29_43 11.551961
Rsp28_44 sp28_44 sp29_44 11.551961
Rsn28_44 sn28_44 sn29_44 11.551961
Rsp28_45 sp28_45 sp29_45 11.551961
Rsn28_45 sn28_45 sn29_45 11.551961
Rsp28_46 sp28_46 sp29_46 11.551961
Rsn28_46 sn28_46 sn29_46 11.551961
Rsp28_47 sp28_47 sp29_47 11.551961
Rsn28_47 sn28_47 sn29_47 11.551961
Rsp28_48 sp28_48 sp29_48 11.551961
Rsn28_48 sn28_48 sn29_48 11.551961
Rsp28_49 sp28_49 sp29_49 11.551961
Rsn28_49 sn28_49 sn29_49 11.551961
Rsp28_50 sp28_50 sp29_50 11.551961
Rsn28_50 sn28_50 sn29_50 11.551961
Rsp28_51 sp28_51 sp29_51 11.551961
Rsn28_51 sn28_51 sn29_51 11.551961
Rsp28_52 sp28_52 sp29_52 11.551961
Rsn28_52 sn28_52 sn29_52 11.551961
Rsp28_53 sp28_53 sp29_53 11.551961
Rsn28_53 sn28_53 sn29_53 11.551961
Rsp28_54 sp28_54 sp29_54 11.551961
Rsn28_54 sn28_54 sn29_54 11.551961
Rsp28_55 sp28_55 sp29_55 11.551961
Rsn28_55 sn28_55 sn29_55 11.551961
Rsp28_56 sp28_56 sp29_56 11.551961
Rsn28_56 sn28_56 sn29_56 11.551961
Rsp28_57 sp28_57 sp29_57 11.551961
Rsn28_57 sn28_57 sn29_57 11.551961
Rsp28_58 sp28_58 sp29_58 11.551961
Rsn28_58 sn28_58 sn29_58 11.551961
Rsp28_59 sp28_59 sp29_59 11.551961
Rsn28_59 sn28_59 sn29_59 11.551961
Rsp28_60 sp28_60 sp29_60 11.551961
Rsn28_60 sn28_60 sn29_60 11.551961
Rsp28_61 sp28_61 sp29_61 11.551961
Rsn28_61 sn28_61 sn29_61 11.551961
Rsp28_62 sp28_62 sp29_62 11.551961
Rsn28_62 sn28_62 sn29_62 11.551961
Rsp28_63 sp28_63 sp29_63 11.551961
Rsn28_63 sn28_63 sn29_63 11.551961
Rsp28_64 sp28_64 sp29_64 11.551961
Rsn28_64 sn28_64 sn29_64 11.551961
Rsp28_65 sp28_65 sp29_65 11.551961
Rsn28_65 sn28_65 sn29_65 11.551961
Rsp28_66 sp28_66 sp29_66 11.551961
Rsn28_66 sn28_66 sn29_66 11.551961
Rsp28_67 sp28_67 sp29_67 11.551961
Rsn28_67 sn28_67 sn29_67 11.551961
Rsp28_68 sp28_68 sp29_68 11.551961
Rsn28_68 sn28_68 sn29_68 11.551961
Rsp28_69 sp28_69 sp29_69 11.551961
Rsn28_69 sn28_69 sn29_69 11.551961
Rsp28_70 sp28_70 sp29_70 11.551961
Rsn28_70 sn28_70 sn29_70 11.551961
Rsp28_71 sp28_71 sp29_71 11.551961
Rsn28_71 sn28_71 sn29_71 11.551961
Rsp28_72 sp28_72 sp29_72 11.551961
Rsn28_72 sn28_72 sn29_72 11.551961
Rsp28_73 sp28_73 sp29_73 11.551961
Rsn28_73 sn28_73 sn29_73 11.551961
Rsp28_74 sp28_74 sp29_74 11.551961
Rsn28_74 sn28_74 sn29_74 11.551961
Rsp28_75 sp28_75 sp29_75 11.551961
Rsn28_75 sn28_75 sn29_75 11.551961
Rsp28_76 sp28_76 sp29_76 11.551961
Rsn28_76 sn28_76 sn29_76 11.551961
Rsp28_77 sp28_77 sp29_77 11.551961
Rsn28_77 sn28_77 sn29_77 11.551961
Rsp28_78 sp28_78 sp29_78 11.551961
Rsn28_78 sn28_78 sn29_78 11.551961
Rsp28_79 sp28_79 sp29_79 11.551961
Rsn28_79 sn28_79 sn29_79 11.551961
Rsp28_80 sp28_80 sp29_80 11.551961
Rsn28_80 sn28_80 sn29_80 11.551961
Rsp28_81 sp28_81 sp29_81 11.551961
Rsn28_81 sn28_81 sn29_81 11.551961
Rsp28_82 sp28_82 sp29_82 11.551961
Rsn28_82 sn28_82 sn29_82 11.551961
Rsp28_83 sp28_83 sp29_83 11.551961
Rsn28_83 sn28_83 sn29_83 11.551961
Rsp28_84 sp28_84 sp29_84 11.551961
Rsn28_84 sn28_84 sn29_84 11.551961
Rsp29_1 sp29_1 sp30_1 11.551961
Rsn29_1 sn29_1 sn30_1 11.551961
Rsp29_2 sp29_2 sp30_2 11.551961
Rsn29_2 sn29_2 sn30_2 11.551961
Rsp29_3 sp29_3 sp30_3 11.551961
Rsn29_3 sn29_3 sn30_3 11.551961
Rsp29_4 sp29_4 sp30_4 11.551961
Rsn29_4 sn29_4 sn30_4 11.551961
Rsp29_5 sp29_5 sp30_5 11.551961
Rsn29_5 sn29_5 sn30_5 11.551961
Rsp29_6 sp29_6 sp30_6 11.551961
Rsn29_6 sn29_6 sn30_6 11.551961
Rsp29_7 sp29_7 sp30_7 11.551961
Rsn29_7 sn29_7 sn30_7 11.551961
Rsp29_8 sp29_8 sp30_8 11.551961
Rsn29_8 sn29_8 sn30_8 11.551961
Rsp29_9 sp29_9 sp30_9 11.551961
Rsn29_9 sn29_9 sn30_9 11.551961
Rsp29_10 sp29_10 sp30_10 11.551961
Rsn29_10 sn29_10 sn30_10 11.551961
Rsp29_11 sp29_11 sp30_11 11.551961
Rsn29_11 sn29_11 sn30_11 11.551961
Rsp29_12 sp29_12 sp30_12 11.551961
Rsn29_12 sn29_12 sn30_12 11.551961
Rsp29_13 sp29_13 sp30_13 11.551961
Rsn29_13 sn29_13 sn30_13 11.551961
Rsp29_14 sp29_14 sp30_14 11.551961
Rsn29_14 sn29_14 sn30_14 11.551961
Rsp29_15 sp29_15 sp30_15 11.551961
Rsn29_15 sn29_15 sn30_15 11.551961
Rsp29_16 sp29_16 sp30_16 11.551961
Rsn29_16 sn29_16 sn30_16 11.551961
Rsp29_17 sp29_17 sp30_17 11.551961
Rsn29_17 sn29_17 sn30_17 11.551961
Rsp29_18 sp29_18 sp30_18 11.551961
Rsn29_18 sn29_18 sn30_18 11.551961
Rsp29_19 sp29_19 sp30_19 11.551961
Rsn29_19 sn29_19 sn30_19 11.551961
Rsp29_20 sp29_20 sp30_20 11.551961
Rsn29_20 sn29_20 sn30_20 11.551961
Rsp29_21 sp29_21 sp30_21 11.551961
Rsn29_21 sn29_21 sn30_21 11.551961
Rsp29_22 sp29_22 sp30_22 11.551961
Rsn29_22 sn29_22 sn30_22 11.551961
Rsp29_23 sp29_23 sp30_23 11.551961
Rsn29_23 sn29_23 sn30_23 11.551961
Rsp29_24 sp29_24 sp30_24 11.551961
Rsn29_24 sn29_24 sn30_24 11.551961
Rsp29_25 sp29_25 sp30_25 11.551961
Rsn29_25 sn29_25 sn30_25 11.551961
Rsp29_26 sp29_26 sp30_26 11.551961
Rsn29_26 sn29_26 sn30_26 11.551961
Rsp29_27 sp29_27 sp30_27 11.551961
Rsn29_27 sn29_27 sn30_27 11.551961
Rsp29_28 sp29_28 sp30_28 11.551961
Rsn29_28 sn29_28 sn30_28 11.551961
Rsp29_29 sp29_29 sp30_29 11.551961
Rsn29_29 sn29_29 sn30_29 11.551961
Rsp29_30 sp29_30 sp30_30 11.551961
Rsn29_30 sn29_30 sn30_30 11.551961
Rsp29_31 sp29_31 sp30_31 11.551961
Rsn29_31 sn29_31 sn30_31 11.551961
Rsp29_32 sp29_32 sp30_32 11.551961
Rsn29_32 sn29_32 sn30_32 11.551961
Rsp29_33 sp29_33 sp30_33 11.551961
Rsn29_33 sn29_33 sn30_33 11.551961
Rsp29_34 sp29_34 sp30_34 11.551961
Rsn29_34 sn29_34 sn30_34 11.551961
Rsp29_35 sp29_35 sp30_35 11.551961
Rsn29_35 sn29_35 sn30_35 11.551961
Rsp29_36 sp29_36 sp30_36 11.551961
Rsn29_36 sn29_36 sn30_36 11.551961
Rsp29_37 sp29_37 sp30_37 11.551961
Rsn29_37 sn29_37 sn30_37 11.551961
Rsp29_38 sp29_38 sp30_38 11.551961
Rsn29_38 sn29_38 sn30_38 11.551961
Rsp29_39 sp29_39 sp30_39 11.551961
Rsn29_39 sn29_39 sn30_39 11.551961
Rsp29_40 sp29_40 sp30_40 11.551961
Rsn29_40 sn29_40 sn30_40 11.551961
Rsp29_41 sp29_41 sp30_41 11.551961
Rsn29_41 sn29_41 sn30_41 11.551961
Rsp29_42 sp29_42 sp30_42 11.551961
Rsn29_42 sn29_42 sn30_42 11.551961
Rsp29_43 sp29_43 sp30_43 11.551961
Rsn29_43 sn29_43 sn30_43 11.551961
Rsp29_44 sp29_44 sp30_44 11.551961
Rsn29_44 sn29_44 sn30_44 11.551961
Rsp29_45 sp29_45 sp30_45 11.551961
Rsn29_45 sn29_45 sn30_45 11.551961
Rsp29_46 sp29_46 sp30_46 11.551961
Rsn29_46 sn29_46 sn30_46 11.551961
Rsp29_47 sp29_47 sp30_47 11.551961
Rsn29_47 sn29_47 sn30_47 11.551961
Rsp29_48 sp29_48 sp30_48 11.551961
Rsn29_48 sn29_48 sn30_48 11.551961
Rsp29_49 sp29_49 sp30_49 11.551961
Rsn29_49 sn29_49 sn30_49 11.551961
Rsp29_50 sp29_50 sp30_50 11.551961
Rsn29_50 sn29_50 sn30_50 11.551961
Rsp29_51 sp29_51 sp30_51 11.551961
Rsn29_51 sn29_51 sn30_51 11.551961
Rsp29_52 sp29_52 sp30_52 11.551961
Rsn29_52 sn29_52 sn30_52 11.551961
Rsp29_53 sp29_53 sp30_53 11.551961
Rsn29_53 sn29_53 sn30_53 11.551961
Rsp29_54 sp29_54 sp30_54 11.551961
Rsn29_54 sn29_54 sn30_54 11.551961
Rsp29_55 sp29_55 sp30_55 11.551961
Rsn29_55 sn29_55 sn30_55 11.551961
Rsp29_56 sp29_56 sp30_56 11.551961
Rsn29_56 sn29_56 sn30_56 11.551961
Rsp29_57 sp29_57 sp30_57 11.551961
Rsn29_57 sn29_57 sn30_57 11.551961
Rsp29_58 sp29_58 sp30_58 11.551961
Rsn29_58 sn29_58 sn30_58 11.551961
Rsp29_59 sp29_59 sp30_59 11.551961
Rsn29_59 sn29_59 sn30_59 11.551961
Rsp29_60 sp29_60 sp30_60 11.551961
Rsn29_60 sn29_60 sn30_60 11.551961
Rsp29_61 sp29_61 sp30_61 11.551961
Rsn29_61 sn29_61 sn30_61 11.551961
Rsp29_62 sp29_62 sp30_62 11.551961
Rsn29_62 sn29_62 sn30_62 11.551961
Rsp29_63 sp29_63 sp30_63 11.551961
Rsn29_63 sn29_63 sn30_63 11.551961
Rsp29_64 sp29_64 sp30_64 11.551961
Rsn29_64 sn29_64 sn30_64 11.551961
Rsp29_65 sp29_65 sp30_65 11.551961
Rsn29_65 sn29_65 sn30_65 11.551961
Rsp29_66 sp29_66 sp30_66 11.551961
Rsn29_66 sn29_66 sn30_66 11.551961
Rsp29_67 sp29_67 sp30_67 11.551961
Rsn29_67 sn29_67 sn30_67 11.551961
Rsp29_68 sp29_68 sp30_68 11.551961
Rsn29_68 sn29_68 sn30_68 11.551961
Rsp29_69 sp29_69 sp30_69 11.551961
Rsn29_69 sn29_69 sn30_69 11.551961
Rsp29_70 sp29_70 sp30_70 11.551961
Rsn29_70 sn29_70 sn30_70 11.551961
Rsp29_71 sp29_71 sp30_71 11.551961
Rsn29_71 sn29_71 sn30_71 11.551961
Rsp29_72 sp29_72 sp30_72 11.551961
Rsn29_72 sn29_72 sn30_72 11.551961
Rsp29_73 sp29_73 sp30_73 11.551961
Rsn29_73 sn29_73 sn30_73 11.551961
Rsp29_74 sp29_74 sp30_74 11.551961
Rsn29_74 sn29_74 sn30_74 11.551961
Rsp29_75 sp29_75 sp30_75 11.551961
Rsn29_75 sn29_75 sn30_75 11.551961
Rsp29_76 sp29_76 sp30_76 11.551961
Rsn29_76 sn29_76 sn30_76 11.551961
Rsp29_77 sp29_77 sp30_77 11.551961
Rsn29_77 sn29_77 sn30_77 11.551961
Rsp29_78 sp29_78 sp30_78 11.551961
Rsn29_78 sn29_78 sn30_78 11.551961
Rsp29_79 sp29_79 sp30_79 11.551961
Rsn29_79 sn29_79 sn30_79 11.551961
Rsp29_80 sp29_80 sp30_80 11.551961
Rsn29_80 sn29_80 sn30_80 11.551961
Rsp29_81 sp29_81 sp30_81 11.551961
Rsn29_81 sn29_81 sn30_81 11.551961
Rsp29_82 sp29_82 sp30_82 11.551961
Rsn29_82 sn29_82 sn30_82 11.551961
Rsp29_83 sp29_83 sp30_83 11.551961
Rsn29_83 sn29_83 sn30_83 11.551961
Rsp29_84 sp29_84 sp30_84 11.551961
Rsn29_84 sn29_84 sn30_84 11.551961
Rsp30_1 sp30_1 sp31_1 11.551961
Rsn30_1 sn30_1 sn31_1 11.551961
Rsp30_2 sp30_2 sp31_2 11.551961
Rsn30_2 sn30_2 sn31_2 11.551961
Rsp30_3 sp30_3 sp31_3 11.551961
Rsn30_3 sn30_3 sn31_3 11.551961
Rsp30_4 sp30_4 sp31_4 11.551961
Rsn30_4 sn30_4 sn31_4 11.551961
Rsp30_5 sp30_5 sp31_5 11.551961
Rsn30_5 sn30_5 sn31_5 11.551961
Rsp30_6 sp30_6 sp31_6 11.551961
Rsn30_6 sn30_6 sn31_6 11.551961
Rsp30_7 sp30_7 sp31_7 11.551961
Rsn30_7 sn30_7 sn31_7 11.551961
Rsp30_8 sp30_8 sp31_8 11.551961
Rsn30_8 sn30_8 sn31_8 11.551961
Rsp30_9 sp30_9 sp31_9 11.551961
Rsn30_9 sn30_9 sn31_9 11.551961
Rsp30_10 sp30_10 sp31_10 11.551961
Rsn30_10 sn30_10 sn31_10 11.551961
Rsp30_11 sp30_11 sp31_11 11.551961
Rsn30_11 sn30_11 sn31_11 11.551961
Rsp30_12 sp30_12 sp31_12 11.551961
Rsn30_12 sn30_12 sn31_12 11.551961
Rsp30_13 sp30_13 sp31_13 11.551961
Rsn30_13 sn30_13 sn31_13 11.551961
Rsp30_14 sp30_14 sp31_14 11.551961
Rsn30_14 sn30_14 sn31_14 11.551961
Rsp30_15 sp30_15 sp31_15 11.551961
Rsn30_15 sn30_15 sn31_15 11.551961
Rsp30_16 sp30_16 sp31_16 11.551961
Rsn30_16 sn30_16 sn31_16 11.551961
Rsp30_17 sp30_17 sp31_17 11.551961
Rsn30_17 sn30_17 sn31_17 11.551961
Rsp30_18 sp30_18 sp31_18 11.551961
Rsn30_18 sn30_18 sn31_18 11.551961
Rsp30_19 sp30_19 sp31_19 11.551961
Rsn30_19 sn30_19 sn31_19 11.551961
Rsp30_20 sp30_20 sp31_20 11.551961
Rsn30_20 sn30_20 sn31_20 11.551961
Rsp30_21 sp30_21 sp31_21 11.551961
Rsn30_21 sn30_21 sn31_21 11.551961
Rsp30_22 sp30_22 sp31_22 11.551961
Rsn30_22 sn30_22 sn31_22 11.551961
Rsp30_23 sp30_23 sp31_23 11.551961
Rsn30_23 sn30_23 sn31_23 11.551961
Rsp30_24 sp30_24 sp31_24 11.551961
Rsn30_24 sn30_24 sn31_24 11.551961
Rsp30_25 sp30_25 sp31_25 11.551961
Rsn30_25 sn30_25 sn31_25 11.551961
Rsp30_26 sp30_26 sp31_26 11.551961
Rsn30_26 sn30_26 sn31_26 11.551961
Rsp30_27 sp30_27 sp31_27 11.551961
Rsn30_27 sn30_27 sn31_27 11.551961
Rsp30_28 sp30_28 sp31_28 11.551961
Rsn30_28 sn30_28 sn31_28 11.551961
Rsp30_29 sp30_29 sp31_29 11.551961
Rsn30_29 sn30_29 sn31_29 11.551961
Rsp30_30 sp30_30 sp31_30 11.551961
Rsn30_30 sn30_30 sn31_30 11.551961
Rsp30_31 sp30_31 sp31_31 11.551961
Rsn30_31 sn30_31 sn31_31 11.551961
Rsp30_32 sp30_32 sp31_32 11.551961
Rsn30_32 sn30_32 sn31_32 11.551961
Rsp30_33 sp30_33 sp31_33 11.551961
Rsn30_33 sn30_33 sn31_33 11.551961
Rsp30_34 sp30_34 sp31_34 11.551961
Rsn30_34 sn30_34 sn31_34 11.551961
Rsp30_35 sp30_35 sp31_35 11.551961
Rsn30_35 sn30_35 sn31_35 11.551961
Rsp30_36 sp30_36 sp31_36 11.551961
Rsn30_36 sn30_36 sn31_36 11.551961
Rsp30_37 sp30_37 sp31_37 11.551961
Rsn30_37 sn30_37 sn31_37 11.551961
Rsp30_38 sp30_38 sp31_38 11.551961
Rsn30_38 sn30_38 sn31_38 11.551961
Rsp30_39 sp30_39 sp31_39 11.551961
Rsn30_39 sn30_39 sn31_39 11.551961
Rsp30_40 sp30_40 sp31_40 11.551961
Rsn30_40 sn30_40 sn31_40 11.551961
Rsp30_41 sp30_41 sp31_41 11.551961
Rsn30_41 sn30_41 sn31_41 11.551961
Rsp30_42 sp30_42 sp31_42 11.551961
Rsn30_42 sn30_42 sn31_42 11.551961
Rsp30_43 sp30_43 sp31_43 11.551961
Rsn30_43 sn30_43 sn31_43 11.551961
Rsp30_44 sp30_44 sp31_44 11.551961
Rsn30_44 sn30_44 sn31_44 11.551961
Rsp30_45 sp30_45 sp31_45 11.551961
Rsn30_45 sn30_45 sn31_45 11.551961
Rsp30_46 sp30_46 sp31_46 11.551961
Rsn30_46 sn30_46 sn31_46 11.551961
Rsp30_47 sp30_47 sp31_47 11.551961
Rsn30_47 sn30_47 sn31_47 11.551961
Rsp30_48 sp30_48 sp31_48 11.551961
Rsn30_48 sn30_48 sn31_48 11.551961
Rsp30_49 sp30_49 sp31_49 11.551961
Rsn30_49 sn30_49 sn31_49 11.551961
Rsp30_50 sp30_50 sp31_50 11.551961
Rsn30_50 sn30_50 sn31_50 11.551961
Rsp30_51 sp30_51 sp31_51 11.551961
Rsn30_51 sn30_51 sn31_51 11.551961
Rsp30_52 sp30_52 sp31_52 11.551961
Rsn30_52 sn30_52 sn31_52 11.551961
Rsp30_53 sp30_53 sp31_53 11.551961
Rsn30_53 sn30_53 sn31_53 11.551961
Rsp30_54 sp30_54 sp31_54 11.551961
Rsn30_54 sn30_54 sn31_54 11.551961
Rsp30_55 sp30_55 sp31_55 11.551961
Rsn30_55 sn30_55 sn31_55 11.551961
Rsp30_56 sp30_56 sp31_56 11.551961
Rsn30_56 sn30_56 sn31_56 11.551961
Rsp30_57 sp30_57 sp31_57 11.551961
Rsn30_57 sn30_57 sn31_57 11.551961
Rsp30_58 sp30_58 sp31_58 11.551961
Rsn30_58 sn30_58 sn31_58 11.551961
Rsp30_59 sp30_59 sp31_59 11.551961
Rsn30_59 sn30_59 sn31_59 11.551961
Rsp30_60 sp30_60 sp31_60 11.551961
Rsn30_60 sn30_60 sn31_60 11.551961
Rsp30_61 sp30_61 sp31_61 11.551961
Rsn30_61 sn30_61 sn31_61 11.551961
Rsp30_62 sp30_62 sp31_62 11.551961
Rsn30_62 sn30_62 sn31_62 11.551961
Rsp30_63 sp30_63 sp31_63 11.551961
Rsn30_63 sn30_63 sn31_63 11.551961
Rsp30_64 sp30_64 sp31_64 11.551961
Rsn30_64 sn30_64 sn31_64 11.551961
Rsp30_65 sp30_65 sp31_65 11.551961
Rsn30_65 sn30_65 sn31_65 11.551961
Rsp30_66 sp30_66 sp31_66 11.551961
Rsn30_66 sn30_66 sn31_66 11.551961
Rsp30_67 sp30_67 sp31_67 11.551961
Rsn30_67 sn30_67 sn31_67 11.551961
Rsp30_68 sp30_68 sp31_68 11.551961
Rsn30_68 sn30_68 sn31_68 11.551961
Rsp30_69 sp30_69 sp31_69 11.551961
Rsn30_69 sn30_69 sn31_69 11.551961
Rsp30_70 sp30_70 sp31_70 11.551961
Rsn30_70 sn30_70 sn31_70 11.551961
Rsp30_71 sp30_71 sp31_71 11.551961
Rsn30_71 sn30_71 sn31_71 11.551961
Rsp30_72 sp30_72 sp31_72 11.551961
Rsn30_72 sn30_72 sn31_72 11.551961
Rsp30_73 sp30_73 sp31_73 11.551961
Rsn30_73 sn30_73 sn31_73 11.551961
Rsp30_74 sp30_74 sp31_74 11.551961
Rsn30_74 sn30_74 sn31_74 11.551961
Rsp30_75 sp30_75 sp31_75 11.551961
Rsn30_75 sn30_75 sn31_75 11.551961
Rsp30_76 sp30_76 sp31_76 11.551961
Rsn30_76 sn30_76 sn31_76 11.551961
Rsp30_77 sp30_77 sp31_77 11.551961
Rsn30_77 sn30_77 sn31_77 11.551961
Rsp30_78 sp30_78 sp31_78 11.551961
Rsn30_78 sn30_78 sn31_78 11.551961
Rsp30_79 sp30_79 sp31_79 11.551961
Rsn30_79 sn30_79 sn31_79 11.551961
Rsp30_80 sp30_80 sp31_80 11.551961
Rsn30_80 sn30_80 sn31_80 11.551961
Rsp30_81 sp30_81 sp31_81 11.551961
Rsn30_81 sn30_81 sn31_81 11.551961
Rsp30_82 sp30_82 sp31_82 11.551961
Rsn30_82 sn30_82 sn31_82 11.551961
Rsp30_83 sp30_83 sp31_83 11.551961
Rsn30_83 sn30_83 sn31_83 11.551961
Rsp30_84 sp30_84 sp31_84 11.551961
Rsn30_84 sn30_84 sn31_84 11.551961
Rsp31_1 sp31_1 sp1_p1 11.551961
Rsn31_1 sn31_1 sn1_p1 11.551961
Rsp31_2 sp31_2 sp2_p1 11.551961
Rsn31_2 sn31_2 sn2_p1 11.551961
Rsp31_3 sp31_3 sp3_p1 11.551961
Rsn31_3 sn31_3 sn3_p1 11.551961
Rsp31_4 sp31_4 sp4_p1 11.551961
Rsn31_4 sn31_4 sn4_p1 11.551961
Rsp31_5 sp31_5 sp5_p1 11.551961
Rsn31_5 sn31_5 sn5_p1 11.551961
Rsp31_6 sp31_6 sp6_p1 11.551961
Rsn31_6 sn31_6 sn6_p1 11.551961
Rsp31_7 sp31_7 sp7_p1 11.551961
Rsn31_7 sn31_7 sn7_p1 11.551961
Rsp31_8 sp31_8 sp8_p1 11.551961
Rsn31_8 sn31_8 sn8_p1 11.551961
Rsp31_9 sp31_9 sp9_p1 11.551961
Rsn31_9 sn31_9 sn9_p1 11.551961
Rsp31_10 sp31_10 sp10_p1 11.551961
Rsn31_10 sn31_10 sn10_p1 11.551961
Rsp31_11 sp31_11 sp11_p1 11.551961
Rsn31_11 sn31_11 sn11_p1 11.551961
Rsp31_12 sp31_12 sp12_p1 11.551961
Rsn31_12 sn31_12 sn12_p1 11.551961
Rsp31_13 sp31_13 sp13_p1 11.551961
Rsn31_13 sn31_13 sn13_p1 11.551961
Rsp31_14 sp31_14 sp14_p1 11.551961
Rsn31_14 sn31_14 sn14_p1 11.551961
Rsp31_15 sp31_15 sp15_p1 11.551961
Rsn31_15 sn31_15 sn15_p1 11.551961
Rsp31_16 sp31_16 sp16_p1 11.551961
Rsn31_16 sn31_16 sn16_p1 11.551961
Rsp31_17 sp31_17 sp17_p1 11.551961
Rsn31_17 sn31_17 sn17_p1 11.551961
Rsp31_18 sp31_18 sp18_p1 11.551961
Rsn31_18 sn31_18 sn18_p1 11.551961
Rsp31_19 sp31_19 sp19_p1 11.551961
Rsn31_19 sn31_19 sn19_p1 11.551961
Rsp31_20 sp31_20 sp20_p1 11.551961
Rsn31_20 sn31_20 sn20_p1 11.551961
Rsp31_21 sp31_21 sp21_p1 11.551961
Rsn31_21 sn31_21 sn21_p1 11.551961
Rsp31_22 sp31_22 sp22_p1 11.551961
Rsn31_22 sn31_22 sn22_p1 11.551961
Rsp31_23 sp31_23 sp23_p1 11.551961
Rsn31_23 sn31_23 sn23_p1 11.551961
Rsp31_24 sp31_24 sp24_p1 11.551961
Rsn31_24 sn31_24 sn24_p1 11.551961
Rsp31_25 sp31_25 sp25_p1 11.551961
Rsn31_25 sn31_25 sn25_p1 11.551961
Rsp31_26 sp31_26 sp26_p1 11.551961
Rsn31_26 sn31_26 sn26_p1 11.551961
Rsp31_27 sp31_27 sp27_p1 11.551961
Rsn31_27 sn31_27 sn27_p1 11.551961
Rsp31_28 sp31_28 sp28_p1 11.551961
Rsn31_28 sn31_28 sn28_p1 11.551961
Rsp31_29 sp31_29 sp29_p1 11.551961
Rsn31_29 sn31_29 sn29_p1 11.551961
Rsp31_30 sp31_30 sp30_p1 11.551961
Rsn31_30 sn31_30 sn30_p1 11.551961
Rsp31_31 sp31_31 sp31_p1 11.551961
Rsn31_31 sn31_31 sn31_p1 11.551961
Rsp31_32 sp31_32 sp32_p1 11.551961
Rsn31_32 sn31_32 sn32_p1 11.551961
Rsp31_33 sp31_33 sp33_p1 11.551961
Rsn31_33 sn31_33 sn33_p1 11.551961
Rsp31_34 sp31_34 sp34_p1 11.551961
Rsn31_34 sn31_34 sn34_p1 11.551961
Rsp31_35 sp31_35 sp35_p1 11.551961
Rsn31_35 sn31_35 sn35_p1 11.551961
Rsp31_36 sp31_36 sp36_p1 11.551961
Rsn31_36 sn31_36 sn36_p1 11.551961
Rsp31_37 sp31_37 sp37_p1 11.551961
Rsn31_37 sn31_37 sn37_p1 11.551961
Rsp31_38 sp31_38 sp38_p1 11.551961
Rsn31_38 sn31_38 sn38_p1 11.551961
Rsp31_39 sp31_39 sp39_p1 11.551961
Rsn31_39 sn31_39 sn39_p1 11.551961
Rsp31_40 sp31_40 sp40_p1 11.551961
Rsn31_40 sn31_40 sn40_p1 11.551961
Rsp31_41 sp31_41 sp41_p1 11.551961
Rsn31_41 sn31_41 sn41_p1 11.551961
Rsp31_42 sp31_42 sp42_p1 11.551961
Rsn31_42 sn31_42 sn42_p1 11.551961
Rsp31_43 sp31_43 sp43_p1 11.551961
Rsn31_43 sn31_43 sn43_p1 11.551961
Rsp31_44 sp31_44 sp44_p1 11.551961
Rsn31_44 sn31_44 sn44_p1 11.551961
Rsp31_45 sp31_45 sp45_p1 11.551961
Rsn31_45 sn31_45 sn45_p1 11.551961
Rsp31_46 sp31_46 sp46_p1 11.551961
Rsn31_46 sn31_46 sn46_p1 11.551961
Rsp31_47 sp31_47 sp47_p1 11.551961
Rsn31_47 sn31_47 sn47_p1 11.551961
Rsp31_48 sp31_48 sp48_p1 11.551961
Rsn31_48 sn31_48 sn48_p1 11.551961
Rsp31_49 sp31_49 sp49_p1 11.551961
Rsn31_49 sn31_49 sn49_p1 11.551961
Rsp31_50 sp31_50 sp50_p1 11.551961
Rsn31_50 sn31_50 sn50_p1 11.551961
Rsp31_51 sp31_51 sp51_p1 11.551961
Rsn31_51 sn31_51 sn51_p1 11.551961
Rsp31_52 sp31_52 sp52_p1 11.551961
Rsn31_52 sn31_52 sn52_p1 11.551961
Rsp31_53 sp31_53 sp53_p1 11.551961
Rsn31_53 sn31_53 sn53_p1 11.551961
Rsp31_54 sp31_54 sp54_p1 11.551961
Rsn31_54 sn31_54 sn54_p1 11.551961
Rsp31_55 sp31_55 sp55_p1 11.551961
Rsn31_55 sn31_55 sn55_p1 11.551961
Rsp31_56 sp31_56 sp56_p1 11.551961
Rsn31_56 sn31_56 sn56_p1 11.551961
Rsp31_57 sp31_57 sp57_p1 11.551961
Rsn31_57 sn31_57 sn57_p1 11.551961
Rsp31_58 sp31_58 sp58_p1 11.551961
Rsn31_58 sn31_58 sn58_p1 11.551961
Rsp31_59 sp31_59 sp59_p1 11.551961
Rsn31_59 sn31_59 sn59_p1 11.551961
Rsp31_60 sp31_60 sp60_p1 11.551961
Rsn31_60 sn31_60 sn60_p1 11.551961
Rsp31_61 sp31_61 sp61_p1 11.551961
Rsn31_61 sn31_61 sn61_p1 11.551961
Rsp31_62 sp31_62 sp62_p1 11.551961
Rsn31_62 sn31_62 sn62_p1 11.551961
Rsp31_63 sp31_63 sp63_p1 11.551961
Rsn31_63 sn31_63 sn63_p1 11.551961
Rsp31_64 sp31_64 sp64_p1 11.551961
Rsn31_64 sn31_64 sn64_p1 11.551961
Rsp31_65 sp31_65 sp65_p1 11.551961
Rsn31_65 sn31_65 sn65_p1 11.551961
Rsp31_66 sp31_66 sp66_p1 11.551961
Rsn31_66 sn31_66 sn66_p1 11.551961
Rsp31_67 sp31_67 sp67_p1 11.551961
Rsn31_67 sn31_67 sn67_p1 11.551961
Rsp31_68 sp31_68 sp68_p1 11.551961
Rsn31_68 sn31_68 sn68_p1 11.551961
Rsp31_69 sp31_69 sp69_p1 11.551961
Rsn31_69 sn31_69 sn69_p1 11.551961
Rsp31_70 sp31_70 sp70_p1 11.551961
Rsn31_70 sn31_70 sn70_p1 11.551961
Rsp31_71 sp31_71 sp71_p1 11.551961
Rsn31_71 sn31_71 sn71_p1 11.551961
Rsp31_72 sp31_72 sp72_p1 11.551961
Rsn31_72 sn31_72 sn72_p1 11.551961
Rsp31_73 sp31_73 sp73_p1 11.551961
Rsn31_73 sn31_73 sn73_p1 11.551961
Rsp31_74 sp31_74 sp74_p1 11.551961
Rsn31_74 sn31_74 sn74_p1 11.551961
Rsp31_75 sp31_75 sp75_p1 11.551961
Rsn31_75 sn31_75 sn75_p1 11.551961
Rsp31_76 sp31_76 sp76_p1 11.551961
Rsn31_76 sn31_76 sn76_p1 11.551961
Rsp31_77 sp31_77 sp77_p1 11.551961
Rsn31_77 sn31_77 sn77_p1 11.551961
Rsp31_78 sp31_78 sp78_p1 11.551961
Rsn31_78 sn31_78 sn78_p1 11.551961
Rsp31_79 sp31_79 sp79_p1 11.551961
Rsn31_79 sn31_79 sn79_p1 11.551961
Rsp31_80 sp31_80 sp80_p1 11.551961
Rsn31_80 sn31_80 sn80_p1 11.551961
Rsp31_81 sp31_81 sp81_p1 11.551961
Rsn31_81 sn31_81 sn81_p1 11.551961
Rsp31_82 sp31_82 sp82_p1 11.551961
Rsn31_82 sn31_82 sn82_p1 11.551961
Rsp31_83 sp31_83 sp83_p1 11.551961
Rsn31_83 sn31_83 sn83_p1 11.551961
Rsp31_84 sp31_84 sp84_p1 11.551961
Rsn31_84 sn31_84 sn84_p1 11.551961
Rsp32_1 sp32_1 sp33_1 11.551961
Rsn32_1 sn32_1 sn33_1 11.551961
Rsp32_2 sp32_2 sp33_2 11.551961
Rsn32_2 sn32_2 sn33_2 11.551961
Rsp32_3 sp32_3 sp33_3 11.551961
Rsn32_3 sn32_3 sn33_3 11.551961
Rsp32_4 sp32_4 sp33_4 11.551961
Rsn32_4 sn32_4 sn33_4 11.551961
Rsp32_5 sp32_5 sp33_5 11.551961
Rsn32_5 sn32_5 sn33_5 11.551961
Rsp32_6 sp32_6 sp33_6 11.551961
Rsn32_6 sn32_6 sn33_6 11.551961
Rsp32_7 sp32_7 sp33_7 11.551961
Rsn32_7 sn32_7 sn33_7 11.551961
Rsp32_8 sp32_8 sp33_8 11.551961
Rsn32_8 sn32_8 sn33_8 11.551961
Rsp32_9 sp32_9 sp33_9 11.551961
Rsn32_9 sn32_9 sn33_9 11.551961
Rsp32_10 sp32_10 sp33_10 11.551961
Rsn32_10 sn32_10 sn33_10 11.551961
Rsp32_11 sp32_11 sp33_11 11.551961
Rsn32_11 sn32_11 sn33_11 11.551961
Rsp32_12 sp32_12 sp33_12 11.551961
Rsn32_12 sn32_12 sn33_12 11.551961
Rsp32_13 sp32_13 sp33_13 11.551961
Rsn32_13 sn32_13 sn33_13 11.551961
Rsp32_14 sp32_14 sp33_14 11.551961
Rsn32_14 sn32_14 sn33_14 11.551961
Rsp32_15 sp32_15 sp33_15 11.551961
Rsn32_15 sn32_15 sn33_15 11.551961
Rsp32_16 sp32_16 sp33_16 11.551961
Rsn32_16 sn32_16 sn33_16 11.551961
Rsp32_17 sp32_17 sp33_17 11.551961
Rsn32_17 sn32_17 sn33_17 11.551961
Rsp32_18 sp32_18 sp33_18 11.551961
Rsn32_18 sn32_18 sn33_18 11.551961
Rsp32_19 sp32_19 sp33_19 11.551961
Rsn32_19 sn32_19 sn33_19 11.551961
Rsp32_20 sp32_20 sp33_20 11.551961
Rsn32_20 sn32_20 sn33_20 11.551961
Rsp32_21 sp32_21 sp33_21 11.551961
Rsn32_21 sn32_21 sn33_21 11.551961
Rsp32_22 sp32_22 sp33_22 11.551961
Rsn32_22 sn32_22 sn33_22 11.551961
Rsp32_23 sp32_23 sp33_23 11.551961
Rsn32_23 sn32_23 sn33_23 11.551961
Rsp32_24 sp32_24 sp33_24 11.551961
Rsn32_24 sn32_24 sn33_24 11.551961
Rsp32_25 sp32_25 sp33_25 11.551961
Rsn32_25 sn32_25 sn33_25 11.551961
Rsp32_26 sp32_26 sp33_26 11.551961
Rsn32_26 sn32_26 sn33_26 11.551961
Rsp32_27 sp32_27 sp33_27 11.551961
Rsn32_27 sn32_27 sn33_27 11.551961
Rsp32_28 sp32_28 sp33_28 11.551961
Rsn32_28 sn32_28 sn33_28 11.551961
Rsp32_29 sp32_29 sp33_29 11.551961
Rsn32_29 sn32_29 sn33_29 11.551961
Rsp32_30 sp32_30 sp33_30 11.551961
Rsn32_30 sn32_30 sn33_30 11.551961
Rsp32_31 sp32_31 sp33_31 11.551961
Rsn32_31 sn32_31 sn33_31 11.551961
Rsp32_32 sp32_32 sp33_32 11.551961
Rsn32_32 sn32_32 sn33_32 11.551961
Rsp32_33 sp32_33 sp33_33 11.551961
Rsn32_33 sn32_33 sn33_33 11.551961
Rsp32_34 sp32_34 sp33_34 11.551961
Rsn32_34 sn32_34 sn33_34 11.551961
Rsp32_35 sp32_35 sp33_35 11.551961
Rsn32_35 sn32_35 sn33_35 11.551961
Rsp32_36 sp32_36 sp33_36 11.551961
Rsn32_36 sn32_36 sn33_36 11.551961
Rsp32_37 sp32_37 sp33_37 11.551961
Rsn32_37 sn32_37 sn33_37 11.551961
Rsp32_38 sp32_38 sp33_38 11.551961
Rsn32_38 sn32_38 sn33_38 11.551961
Rsp32_39 sp32_39 sp33_39 11.551961
Rsn32_39 sn32_39 sn33_39 11.551961
Rsp32_40 sp32_40 sp33_40 11.551961
Rsn32_40 sn32_40 sn33_40 11.551961
Rsp32_41 sp32_41 sp33_41 11.551961
Rsn32_41 sn32_41 sn33_41 11.551961
Rsp32_42 sp32_42 sp33_42 11.551961
Rsn32_42 sn32_42 sn33_42 11.551961
Rsp32_43 sp32_43 sp33_43 11.551961
Rsn32_43 sn32_43 sn33_43 11.551961
Rsp32_44 sp32_44 sp33_44 11.551961
Rsn32_44 sn32_44 sn33_44 11.551961
Rsp32_45 sp32_45 sp33_45 11.551961
Rsn32_45 sn32_45 sn33_45 11.551961
Rsp32_46 sp32_46 sp33_46 11.551961
Rsn32_46 sn32_46 sn33_46 11.551961
Rsp32_47 sp32_47 sp33_47 11.551961
Rsn32_47 sn32_47 sn33_47 11.551961
Rsp32_48 sp32_48 sp33_48 11.551961
Rsn32_48 sn32_48 sn33_48 11.551961
Rsp32_49 sp32_49 sp33_49 11.551961
Rsn32_49 sn32_49 sn33_49 11.551961
Rsp32_50 sp32_50 sp33_50 11.551961
Rsn32_50 sn32_50 sn33_50 11.551961
Rsp32_51 sp32_51 sp33_51 11.551961
Rsn32_51 sn32_51 sn33_51 11.551961
Rsp32_52 sp32_52 sp33_52 11.551961
Rsn32_52 sn32_52 sn33_52 11.551961
Rsp32_53 sp32_53 sp33_53 11.551961
Rsn32_53 sn32_53 sn33_53 11.551961
Rsp32_54 sp32_54 sp33_54 11.551961
Rsn32_54 sn32_54 sn33_54 11.551961
Rsp32_55 sp32_55 sp33_55 11.551961
Rsn32_55 sn32_55 sn33_55 11.551961
Rsp32_56 sp32_56 sp33_56 11.551961
Rsn32_56 sn32_56 sn33_56 11.551961
Rsp32_57 sp32_57 sp33_57 11.551961
Rsn32_57 sn32_57 sn33_57 11.551961
Rsp32_58 sp32_58 sp33_58 11.551961
Rsn32_58 sn32_58 sn33_58 11.551961
Rsp32_59 sp32_59 sp33_59 11.551961
Rsn32_59 sn32_59 sn33_59 11.551961
Rsp32_60 sp32_60 sp33_60 11.551961
Rsn32_60 sn32_60 sn33_60 11.551961
Rsp32_61 sp32_61 sp33_61 11.551961
Rsn32_61 sn32_61 sn33_61 11.551961
Rsp32_62 sp32_62 sp33_62 11.551961
Rsn32_62 sn32_62 sn33_62 11.551961
Rsp32_63 sp32_63 sp33_63 11.551961
Rsn32_63 sn32_63 sn33_63 11.551961
Rsp32_64 sp32_64 sp33_64 11.551961
Rsn32_64 sn32_64 sn33_64 11.551961
Rsp32_65 sp32_65 sp33_65 11.551961
Rsn32_65 sn32_65 sn33_65 11.551961
Rsp32_66 sp32_66 sp33_66 11.551961
Rsn32_66 sn32_66 sn33_66 11.551961
Rsp32_67 sp32_67 sp33_67 11.551961
Rsn32_67 sn32_67 sn33_67 11.551961
Rsp32_68 sp32_68 sp33_68 11.551961
Rsn32_68 sn32_68 sn33_68 11.551961
Rsp32_69 sp32_69 sp33_69 11.551961
Rsn32_69 sn32_69 sn33_69 11.551961
Rsp32_70 sp32_70 sp33_70 11.551961
Rsn32_70 sn32_70 sn33_70 11.551961
Rsp32_71 sp32_71 sp33_71 11.551961
Rsn32_71 sn32_71 sn33_71 11.551961
Rsp32_72 sp32_72 sp33_72 11.551961
Rsn32_72 sn32_72 sn33_72 11.551961
Rsp32_73 sp32_73 sp33_73 11.551961
Rsn32_73 sn32_73 sn33_73 11.551961
Rsp32_74 sp32_74 sp33_74 11.551961
Rsn32_74 sn32_74 sn33_74 11.551961
Rsp32_75 sp32_75 sp33_75 11.551961
Rsn32_75 sn32_75 sn33_75 11.551961
Rsp32_76 sp32_76 sp33_76 11.551961
Rsn32_76 sn32_76 sn33_76 11.551961
Rsp32_77 sp32_77 sp33_77 11.551961
Rsn32_77 sn32_77 sn33_77 11.551961
Rsp32_78 sp32_78 sp33_78 11.551961
Rsn32_78 sn32_78 sn33_78 11.551961
Rsp32_79 sp32_79 sp33_79 11.551961
Rsn32_79 sn32_79 sn33_79 11.551961
Rsp32_80 sp32_80 sp33_80 11.551961
Rsn32_80 sn32_80 sn33_80 11.551961
Rsp32_81 sp32_81 sp33_81 11.551961
Rsn32_81 sn32_81 sn33_81 11.551961
Rsp32_82 sp32_82 sp33_82 11.551961
Rsn32_82 sn32_82 sn33_82 11.551961
Rsp32_83 sp32_83 sp33_83 11.551961
Rsn32_83 sn32_83 sn33_83 11.551961
Rsp32_84 sp32_84 sp33_84 11.551961
Rsn32_84 sn32_84 sn33_84 11.551961
Rsp33_1 sp33_1 sp34_1 11.551961
Rsn33_1 sn33_1 sn34_1 11.551961
Rsp33_2 sp33_2 sp34_2 11.551961
Rsn33_2 sn33_2 sn34_2 11.551961
Rsp33_3 sp33_3 sp34_3 11.551961
Rsn33_3 sn33_3 sn34_3 11.551961
Rsp33_4 sp33_4 sp34_4 11.551961
Rsn33_4 sn33_4 sn34_4 11.551961
Rsp33_5 sp33_5 sp34_5 11.551961
Rsn33_5 sn33_5 sn34_5 11.551961
Rsp33_6 sp33_6 sp34_6 11.551961
Rsn33_6 sn33_6 sn34_6 11.551961
Rsp33_7 sp33_7 sp34_7 11.551961
Rsn33_7 sn33_7 sn34_7 11.551961
Rsp33_8 sp33_8 sp34_8 11.551961
Rsn33_8 sn33_8 sn34_8 11.551961
Rsp33_9 sp33_9 sp34_9 11.551961
Rsn33_9 sn33_9 sn34_9 11.551961
Rsp33_10 sp33_10 sp34_10 11.551961
Rsn33_10 sn33_10 sn34_10 11.551961
Rsp33_11 sp33_11 sp34_11 11.551961
Rsn33_11 sn33_11 sn34_11 11.551961
Rsp33_12 sp33_12 sp34_12 11.551961
Rsn33_12 sn33_12 sn34_12 11.551961
Rsp33_13 sp33_13 sp34_13 11.551961
Rsn33_13 sn33_13 sn34_13 11.551961
Rsp33_14 sp33_14 sp34_14 11.551961
Rsn33_14 sn33_14 sn34_14 11.551961
Rsp33_15 sp33_15 sp34_15 11.551961
Rsn33_15 sn33_15 sn34_15 11.551961
Rsp33_16 sp33_16 sp34_16 11.551961
Rsn33_16 sn33_16 sn34_16 11.551961
Rsp33_17 sp33_17 sp34_17 11.551961
Rsn33_17 sn33_17 sn34_17 11.551961
Rsp33_18 sp33_18 sp34_18 11.551961
Rsn33_18 sn33_18 sn34_18 11.551961
Rsp33_19 sp33_19 sp34_19 11.551961
Rsn33_19 sn33_19 sn34_19 11.551961
Rsp33_20 sp33_20 sp34_20 11.551961
Rsn33_20 sn33_20 sn34_20 11.551961
Rsp33_21 sp33_21 sp34_21 11.551961
Rsn33_21 sn33_21 sn34_21 11.551961
Rsp33_22 sp33_22 sp34_22 11.551961
Rsn33_22 sn33_22 sn34_22 11.551961
Rsp33_23 sp33_23 sp34_23 11.551961
Rsn33_23 sn33_23 sn34_23 11.551961
Rsp33_24 sp33_24 sp34_24 11.551961
Rsn33_24 sn33_24 sn34_24 11.551961
Rsp33_25 sp33_25 sp34_25 11.551961
Rsn33_25 sn33_25 sn34_25 11.551961
Rsp33_26 sp33_26 sp34_26 11.551961
Rsn33_26 sn33_26 sn34_26 11.551961
Rsp33_27 sp33_27 sp34_27 11.551961
Rsn33_27 sn33_27 sn34_27 11.551961
Rsp33_28 sp33_28 sp34_28 11.551961
Rsn33_28 sn33_28 sn34_28 11.551961
Rsp33_29 sp33_29 sp34_29 11.551961
Rsn33_29 sn33_29 sn34_29 11.551961
Rsp33_30 sp33_30 sp34_30 11.551961
Rsn33_30 sn33_30 sn34_30 11.551961
Rsp33_31 sp33_31 sp34_31 11.551961
Rsn33_31 sn33_31 sn34_31 11.551961
Rsp33_32 sp33_32 sp34_32 11.551961
Rsn33_32 sn33_32 sn34_32 11.551961
Rsp33_33 sp33_33 sp34_33 11.551961
Rsn33_33 sn33_33 sn34_33 11.551961
Rsp33_34 sp33_34 sp34_34 11.551961
Rsn33_34 sn33_34 sn34_34 11.551961
Rsp33_35 sp33_35 sp34_35 11.551961
Rsn33_35 sn33_35 sn34_35 11.551961
Rsp33_36 sp33_36 sp34_36 11.551961
Rsn33_36 sn33_36 sn34_36 11.551961
Rsp33_37 sp33_37 sp34_37 11.551961
Rsn33_37 sn33_37 sn34_37 11.551961
Rsp33_38 sp33_38 sp34_38 11.551961
Rsn33_38 sn33_38 sn34_38 11.551961
Rsp33_39 sp33_39 sp34_39 11.551961
Rsn33_39 sn33_39 sn34_39 11.551961
Rsp33_40 sp33_40 sp34_40 11.551961
Rsn33_40 sn33_40 sn34_40 11.551961
Rsp33_41 sp33_41 sp34_41 11.551961
Rsn33_41 sn33_41 sn34_41 11.551961
Rsp33_42 sp33_42 sp34_42 11.551961
Rsn33_42 sn33_42 sn34_42 11.551961
Rsp33_43 sp33_43 sp34_43 11.551961
Rsn33_43 sn33_43 sn34_43 11.551961
Rsp33_44 sp33_44 sp34_44 11.551961
Rsn33_44 sn33_44 sn34_44 11.551961
Rsp33_45 sp33_45 sp34_45 11.551961
Rsn33_45 sn33_45 sn34_45 11.551961
Rsp33_46 sp33_46 sp34_46 11.551961
Rsn33_46 sn33_46 sn34_46 11.551961
Rsp33_47 sp33_47 sp34_47 11.551961
Rsn33_47 sn33_47 sn34_47 11.551961
Rsp33_48 sp33_48 sp34_48 11.551961
Rsn33_48 sn33_48 sn34_48 11.551961
Rsp33_49 sp33_49 sp34_49 11.551961
Rsn33_49 sn33_49 sn34_49 11.551961
Rsp33_50 sp33_50 sp34_50 11.551961
Rsn33_50 sn33_50 sn34_50 11.551961
Rsp33_51 sp33_51 sp34_51 11.551961
Rsn33_51 sn33_51 sn34_51 11.551961
Rsp33_52 sp33_52 sp34_52 11.551961
Rsn33_52 sn33_52 sn34_52 11.551961
Rsp33_53 sp33_53 sp34_53 11.551961
Rsn33_53 sn33_53 sn34_53 11.551961
Rsp33_54 sp33_54 sp34_54 11.551961
Rsn33_54 sn33_54 sn34_54 11.551961
Rsp33_55 sp33_55 sp34_55 11.551961
Rsn33_55 sn33_55 sn34_55 11.551961
Rsp33_56 sp33_56 sp34_56 11.551961
Rsn33_56 sn33_56 sn34_56 11.551961
Rsp33_57 sp33_57 sp34_57 11.551961
Rsn33_57 sn33_57 sn34_57 11.551961
Rsp33_58 sp33_58 sp34_58 11.551961
Rsn33_58 sn33_58 sn34_58 11.551961
Rsp33_59 sp33_59 sp34_59 11.551961
Rsn33_59 sn33_59 sn34_59 11.551961
Rsp33_60 sp33_60 sp34_60 11.551961
Rsn33_60 sn33_60 sn34_60 11.551961
Rsp33_61 sp33_61 sp34_61 11.551961
Rsn33_61 sn33_61 sn34_61 11.551961
Rsp33_62 sp33_62 sp34_62 11.551961
Rsn33_62 sn33_62 sn34_62 11.551961
Rsp33_63 sp33_63 sp34_63 11.551961
Rsn33_63 sn33_63 sn34_63 11.551961
Rsp33_64 sp33_64 sp34_64 11.551961
Rsn33_64 sn33_64 sn34_64 11.551961
Rsp33_65 sp33_65 sp34_65 11.551961
Rsn33_65 sn33_65 sn34_65 11.551961
Rsp33_66 sp33_66 sp34_66 11.551961
Rsn33_66 sn33_66 sn34_66 11.551961
Rsp33_67 sp33_67 sp34_67 11.551961
Rsn33_67 sn33_67 sn34_67 11.551961
Rsp33_68 sp33_68 sp34_68 11.551961
Rsn33_68 sn33_68 sn34_68 11.551961
Rsp33_69 sp33_69 sp34_69 11.551961
Rsn33_69 sn33_69 sn34_69 11.551961
Rsp33_70 sp33_70 sp34_70 11.551961
Rsn33_70 sn33_70 sn34_70 11.551961
Rsp33_71 sp33_71 sp34_71 11.551961
Rsn33_71 sn33_71 sn34_71 11.551961
Rsp33_72 sp33_72 sp34_72 11.551961
Rsn33_72 sn33_72 sn34_72 11.551961
Rsp33_73 sp33_73 sp34_73 11.551961
Rsn33_73 sn33_73 sn34_73 11.551961
Rsp33_74 sp33_74 sp34_74 11.551961
Rsn33_74 sn33_74 sn34_74 11.551961
Rsp33_75 sp33_75 sp34_75 11.551961
Rsn33_75 sn33_75 sn34_75 11.551961
Rsp33_76 sp33_76 sp34_76 11.551961
Rsn33_76 sn33_76 sn34_76 11.551961
Rsp33_77 sp33_77 sp34_77 11.551961
Rsn33_77 sn33_77 sn34_77 11.551961
Rsp33_78 sp33_78 sp34_78 11.551961
Rsn33_78 sn33_78 sn34_78 11.551961
Rsp33_79 sp33_79 sp34_79 11.551961
Rsn33_79 sn33_79 sn34_79 11.551961
Rsp33_80 sp33_80 sp34_80 11.551961
Rsn33_80 sn33_80 sn34_80 11.551961
Rsp33_81 sp33_81 sp34_81 11.551961
Rsn33_81 sn33_81 sn34_81 11.551961
Rsp33_82 sp33_82 sp34_82 11.551961
Rsn33_82 sn33_82 sn34_82 11.551961
Rsp33_83 sp33_83 sp34_83 11.551961
Rsn33_83 sn33_83 sn34_83 11.551961
Rsp33_84 sp33_84 sp34_84 11.551961
Rsn33_84 sn33_84 sn34_84 11.551961
Rsp34_1 sp34_1 sp35_1 11.551961
Rsn34_1 sn34_1 sn35_1 11.551961
Rsp34_2 sp34_2 sp35_2 11.551961
Rsn34_2 sn34_2 sn35_2 11.551961
Rsp34_3 sp34_3 sp35_3 11.551961
Rsn34_3 sn34_3 sn35_3 11.551961
Rsp34_4 sp34_4 sp35_4 11.551961
Rsn34_4 sn34_4 sn35_4 11.551961
Rsp34_5 sp34_5 sp35_5 11.551961
Rsn34_5 sn34_5 sn35_5 11.551961
Rsp34_6 sp34_6 sp35_6 11.551961
Rsn34_6 sn34_6 sn35_6 11.551961
Rsp34_7 sp34_7 sp35_7 11.551961
Rsn34_7 sn34_7 sn35_7 11.551961
Rsp34_8 sp34_8 sp35_8 11.551961
Rsn34_8 sn34_8 sn35_8 11.551961
Rsp34_9 sp34_9 sp35_9 11.551961
Rsn34_9 sn34_9 sn35_9 11.551961
Rsp34_10 sp34_10 sp35_10 11.551961
Rsn34_10 sn34_10 sn35_10 11.551961
Rsp34_11 sp34_11 sp35_11 11.551961
Rsn34_11 sn34_11 sn35_11 11.551961
Rsp34_12 sp34_12 sp35_12 11.551961
Rsn34_12 sn34_12 sn35_12 11.551961
Rsp34_13 sp34_13 sp35_13 11.551961
Rsn34_13 sn34_13 sn35_13 11.551961
Rsp34_14 sp34_14 sp35_14 11.551961
Rsn34_14 sn34_14 sn35_14 11.551961
Rsp34_15 sp34_15 sp35_15 11.551961
Rsn34_15 sn34_15 sn35_15 11.551961
Rsp34_16 sp34_16 sp35_16 11.551961
Rsn34_16 sn34_16 sn35_16 11.551961
Rsp34_17 sp34_17 sp35_17 11.551961
Rsn34_17 sn34_17 sn35_17 11.551961
Rsp34_18 sp34_18 sp35_18 11.551961
Rsn34_18 sn34_18 sn35_18 11.551961
Rsp34_19 sp34_19 sp35_19 11.551961
Rsn34_19 sn34_19 sn35_19 11.551961
Rsp34_20 sp34_20 sp35_20 11.551961
Rsn34_20 sn34_20 sn35_20 11.551961
Rsp34_21 sp34_21 sp35_21 11.551961
Rsn34_21 sn34_21 sn35_21 11.551961
Rsp34_22 sp34_22 sp35_22 11.551961
Rsn34_22 sn34_22 sn35_22 11.551961
Rsp34_23 sp34_23 sp35_23 11.551961
Rsn34_23 sn34_23 sn35_23 11.551961
Rsp34_24 sp34_24 sp35_24 11.551961
Rsn34_24 sn34_24 sn35_24 11.551961
Rsp34_25 sp34_25 sp35_25 11.551961
Rsn34_25 sn34_25 sn35_25 11.551961
Rsp34_26 sp34_26 sp35_26 11.551961
Rsn34_26 sn34_26 sn35_26 11.551961
Rsp34_27 sp34_27 sp35_27 11.551961
Rsn34_27 sn34_27 sn35_27 11.551961
Rsp34_28 sp34_28 sp35_28 11.551961
Rsn34_28 sn34_28 sn35_28 11.551961
Rsp34_29 sp34_29 sp35_29 11.551961
Rsn34_29 sn34_29 sn35_29 11.551961
Rsp34_30 sp34_30 sp35_30 11.551961
Rsn34_30 sn34_30 sn35_30 11.551961
Rsp34_31 sp34_31 sp35_31 11.551961
Rsn34_31 sn34_31 sn35_31 11.551961
Rsp34_32 sp34_32 sp35_32 11.551961
Rsn34_32 sn34_32 sn35_32 11.551961
Rsp34_33 sp34_33 sp35_33 11.551961
Rsn34_33 sn34_33 sn35_33 11.551961
Rsp34_34 sp34_34 sp35_34 11.551961
Rsn34_34 sn34_34 sn35_34 11.551961
Rsp34_35 sp34_35 sp35_35 11.551961
Rsn34_35 sn34_35 sn35_35 11.551961
Rsp34_36 sp34_36 sp35_36 11.551961
Rsn34_36 sn34_36 sn35_36 11.551961
Rsp34_37 sp34_37 sp35_37 11.551961
Rsn34_37 sn34_37 sn35_37 11.551961
Rsp34_38 sp34_38 sp35_38 11.551961
Rsn34_38 sn34_38 sn35_38 11.551961
Rsp34_39 sp34_39 sp35_39 11.551961
Rsn34_39 sn34_39 sn35_39 11.551961
Rsp34_40 sp34_40 sp35_40 11.551961
Rsn34_40 sn34_40 sn35_40 11.551961
Rsp34_41 sp34_41 sp35_41 11.551961
Rsn34_41 sn34_41 sn35_41 11.551961
Rsp34_42 sp34_42 sp35_42 11.551961
Rsn34_42 sn34_42 sn35_42 11.551961
Rsp34_43 sp34_43 sp35_43 11.551961
Rsn34_43 sn34_43 sn35_43 11.551961
Rsp34_44 sp34_44 sp35_44 11.551961
Rsn34_44 sn34_44 sn35_44 11.551961
Rsp34_45 sp34_45 sp35_45 11.551961
Rsn34_45 sn34_45 sn35_45 11.551961
Rsp34_46 sp34_46 sp35_46 11.551961
Rsn34_46 sn34_46 sn35_46 11.551961
Rsp34_47 sp34_47 sp35_47 11.551961
Rsn34_47 sn34_47 sn35_47 11.551961
Rsp34_48 sp34_48 sp35_48 11.551961
Rsn34_48 sn34_48 sn35_48 11.551961
Rsp34_49 sp34_49 sp35_49 11.551961
Rsn34_49 sn34_49 sn35_49 11.551961
Rsp34_50 sp34_50 sp35_50 11.551961
Rsn34_50 sn34_50 sn35_50 11.551961
Rsp34_51 sp34_51 sp35_51 11.551961
Rsn34_51 sn34_51 sn35_51 11.551961
Rsp34_52 sp34_52 sp35_52 11.551961
Rsn34_52 sn34_52 sn35_52 11.551961
Rsp34_53 sp34_53 sp35_53 11.551961
Rsn34_53 sn34_53 sn35_53 11.551961
Rsp34_54 sp34_54 sp35_54 11.551961
Rsn34_54 sn34_54 sn35_54 11.551961
Rsp34_55 sp34_55 sp35_55 11.551961
Rsn34_55 sn34_55 sn35_55 11.551961
Rsp34_56 sp34_56 sp35_56 11.551961
Rsn34_56 sn34_56 sn35_56 11.551961
Rsp34_57 sp34_57 sp35_57 11.551961
Rsn34_57 sn34_57 sn35_57 11.551961
Rsp34_58 sp34_58 sp35_58 11.551961
Rsn34_58 sn34_58 sn35_58 11.551961
Rsp34_59 sp34_59 sp35_59 11.551961
Rsn34_59 sn34_59 sn35_59 11.551961
Rsp34_60 sp34_60 sp35_60 11.551961
Rsn34_60 sn34_60 sn35_60 11.551961
Rsp34_61 sp34_61 sp35_61 11.551961
Rsn34_61 sn34_61 sn35_61 11.551961
Rsp34_62 sp34_62 sp35_62 11.551961
Rsn34_62 sn34_62 sn35_62 11.551961
Rsp34_63 sp34_63 sp35_63 11.551961
Rsn34_63 sn34_63 sn35_63 11.551961
Rsp34_64 sp34_64 sp35_64 11.551961
Rsn34_64 sn34_64 sn35_64 11.551961
Rsp34_65 sp34_65 sp35_65 11.551961
Rsn34_65 sn34_65 sn35_65 11.551961
Rsp34_66 sp34_66 sp35_66 11.551961
Rsn34_66 sn34_66 sn35_66 11.551961
Rsp34_67 sp34_67 sp35_67 11.551961
Rsn34_67 sn34_67 sn35_67 11.551961
Rsp34_68 sp34_68 sp35_68 11.551961
Rsn34_68 sn34_68 sn35_68 11.551961
Rsp34_69 sp34_69 sp35_69 11.551961
Rsn34_69 sn34_69 sn35_69 11.551961
Rsp34_70 sp34_70 sp35_70 11.551961
Rsn34_70 sn34_70 sn35_70 11.551961
Rsp34_71 sp34_71 sp35_71 11.551961
Rsn34_71 sn34_71 sn35_71 11.551961
Rsp34_72 sp34_72 sp35_72 11.551961
Rsn34_72 sn34_72 sn35_72 11.551961
Rsp34_73 sp34_73 sp35_73 11.551961
Rsn34_73 sn34_73 sn35_73 11.551961
Rsp34_74 sp34_74 sp35_74 11.551961
Rsn34_74 sn34_74 sn35_74 11.551961
Rsp34_75 sp34_75 sp35_75 11.551961
Rsn34_75 sn34_75 sn35_75 11.551961
Rsp34_76 sp34_76 sp35_76 11.551961
Rsn34_76 sn34_76 sn35_76 11.551961
Rsp34_77 sp34_77 sp35_77 11.551961
Rsn34_77 sn34_77 sn35_77 11.551961
Rsp34_78 sp34_78 sp35_78 11.551961
Rsn34_78 sn34_78 sn35_78 11.551961
Rsp34_79 sp34_79 sp35_79 11.551961
Rsn34_79 sn34_79 sn35_79 11.551961
Rsp34_80 sp34_80 sp35_80 11.551961
Rsn34_80 sn34_80 sn35_80 11.551961
Rsp34_81 sp34_81 sp35_81 11.551961
Rsn34_81 sn34_81 sn35_81 11.551961
Rsp34_82 sp34_82 sp35_82 11.551961
Rsn34_82 sn34_82 sn35_82 11.551961
Rsp34_83 sp34_83 sp35_83 11.551961
Rsn34_83 sn34_83 sn35_83 11.551961
Rsp34_84 sp34_84 sp35_84 11.551961
Rsn34_84 sn34_84 sn35_84 11.551961
Rsp35_1 sp35_1 sp36_1 11.551961
Rsn35_1 sn35_1 sn36_1 11.551961
Rsp35_2 sp35_2 sp36_2 11.551961
Rsn35_2 sn35_2 sn36_2 11.551961
Rsp35_3 sp35_3 sp36_3 11.551961
Rsn35_3 sn35_3 sn36_3 11.551961
Rsp35_4 sp35_4 sp36_4 11.551961
Rsn35_4 sn35_4 sn36_4 11.551961
Rsp35_5 sp35_5 sp36_5 11.551961
Rsn35_5 sn35_5 sn36_5 11.551961
Rsp35_6 sp35_6 sp36_6 11.551961
Rsn35_6 sn35_6 sn36_6 11.551961
Rsp35_7 sp35_7 sp36_7 11.551961
Rsn35_7 sn35_7 sn36_7 11.551961
Rsp35_8 sp35_8 sp36_8 11.551961
Rsn35_8 sn35_8 sn36_8 11.551961
Rsp35_9 sp35_9 sp36_9 11.551961
Rsn35_9 sn35_9 sn36_9 11.551961
Rsp35_10 sp35_10 sp36_10 11.551961
Rsn35_10 sn35_10 sn36_10 11.551961
Rsp35_11 sp35_11 sp36_11 11.551961
Rsn35_11 sn35_11 sn36_11 11.551961
Rsp35_12 sp35_12 sp36_12 11.551961
Rsn35_12 sn35_12 sn36_12 11.551961
Rsp35_13 sp35_13 sp36_13 11.551961
Rsn35_13 sn35_13 sn36_13 11.551961
Rsp35_14 sp35_14 sp36_14 11.551961
Rsn35_14 sn35_14 sn36_14 11.551961
Rsp35_15 sp35_15 sp36_15 11.551961
Rsn35_15 sn35_15 sn36_15 11.551961
Rsp35_16 sp35_16 sp36_16 11.551961
Rsn35_16 sn35_16 sn36_16 11.551961
Rsp35_17 sp35_17 sp36_17 11.551961
Rsn35_17 sn35_17 sn36_17 11.551961
Rsp35_18 sp35_18 sp36_18 11.551961
Rsn35_18 sn35_18 sn36_18 11.551961
Rsp35_19 sp35_19 sp36_19 11.551961
Rsn35_19 sn35_19 sn36_19 11.551961
Rsp35_20 sp35_20 sp36_20 11.551961
Rsn35_20 sn35_20 sn36_20 11.551961
Rsp35_21 sp35_21 sp36_21 11.551961
Rsn35_21 sn35_21 sn36_21 11.551961
Rsp35_22 sp35_22 sp36_22 11.551961
Rsn35_22 sn35_22 sn36_22 11.551961
Rsp35_23 sp35_23 sp36_23 11.551961
Rsn35_23 sn35_23 sn36_23 11.551961
Rsp35_24 sp35_24 sp36_24 11.551961
Rsn35_24 sn35_24 sn36_24 11.551961
Rsp35_25 sp35_25 sp36_25 11.551961
Rsn35_25 sn35_25 sn36_25 11.551961
Rsp35_26 sp35_26 sp36_26 11.551961
Rsn35_26 sn35_26 sn36_26 11.551961
Rsp35_27 sp35_27 sp36_27 11.551961
Rsn35_27 sn35_27 sn36_27 11.551961
Rsp35_28 sp35_28 sp36_28 11.551961
Rsn35_28 sn35_28 sn36_28 11.551961
Rsp35_29 sp35_29 sp36_29 11.551961
Rsn35_29 sn35_29 sn36_29 11.551961
Rsp35_30 sp35_30 sp36_30 11.551961
Rsn35_30 sn35_30 sn36_30 11.551961
Rsp35_31 sp35_31 sp36_31 11.551961
Rsn35_31 sn35_31 sn36_31 11.551961
Rsp35_32 sp35_32 sp36_32 11.551961
Rsn35_32 sn35_32 sn36_32 11.551961
Rsp35_33 sp35_33 sp36_33 11.551961
Rsn35_33 sn35_33 sn36_33 11.551961
Rsp35_34 sp35_34 sp36_34 11.551961
Rsn35_34 sn35_34 sn36_34 11.551961
Rsp35_35 sp35_35 sp36_35 11.551961
Rsn35_35 sn35_35 sn36_35 11.551961
Rsp35_36 sp35_36 sp36_36 11.551961
Rsn35_36 sn35_36 sn36_36 11.551961
Rsp35_37 sp35_37 sp36_37 11.551961
Rsn35_37 sn35_37 sn36_37 11.551961
Rsp35_38 sp35_38 sp36_38 11.551961
Rsn35_38 sn35_38 sn36_38 11.551961
Rsp35_39 sp35_39 sp36_39 11.551961
Rsn35_39 sn35_39 sn36_39 11.551961
Rsp35_40 sp35_40 sp36_40 11.551961
Rsn35_40 sn35_40 sn36_40 11.551961
Rsp35_41 sp35_41 sp36_41 11.551961
Rsn35_41 sn35_41 sn36_41 11.551961
Rsp35_42 sp35_42 sp36_42 11.551961
Rsn35_42 sn35_42 sn36_42 11.551961
Rsp35_43 sp35_43 sp36_43 11.551961
Rsn35_43 sn35_43 sn36_43 11.551961
Rsp35_44 sp35_44 sp36_44 11.551961
Rsn35_44 sn35_44 sn36_44 11.551961
Rsp35_45 sp35_45 sp36_45 11.551961
Rsn35_45 sn35_45 sn36_45 11.551961
Rsp35_46 sp35_46 sp36_46 11.551961
Rsn35_46 sn35_46 sn36_46 11.551961
Rsp35_47 sp35_47 sp36_47 11.551961
Rsn35_47 sn35_47 sn36_47 11.551961
Rsp35_48 sp35_48 sp36_48 11.551961
Rsn35_48 sn35_48 sn36_48 11.551961
Rsp35_49 sp35_49 sp36_49 11.551961
Rsn35_49 sn35_49 sn36_49 11.551961
Rsp35_50 sp35_50 sp36_50 11.551961
Rsn35_50 sn35_50 sn36_50 11.551961
Rsp35_51 sp35_51 sp36_51 11.551961
Rsn35_51 sn35_51 sn36_51 11.551961
Rsp35_52 sp35_52 sp36_52 11.551961
Rsn35_52 sn35_52 sn36_52 11.551961
Rsp35_53 sp35_53 sp36_53 11.551961
Rsn35_53 sn35_53 sn36_53 11.551961
Rsp35_54 sp35_54 sp36_54 11.551961
Rsn35_54 sn35_54 sn36_54 11.551961
Rsp35_55 sp35_55 sp36_55 11.551961
Rsn35_55 sn35_55 sn36_55 11.551961
Rsp35_56 sp35_56 sp36_56 11.551961
Rsn35_56 sn35_56 sn36_56 11.551961
Rsp35_57 sp35_57 sp36_57 11.551961
Rsn35_57 sn35_57 sn36_57 11.551961
Rsp35_58 sp35_58 sp36_58 11.551961
Rsn35_58 sn35_58 sn36_58 11.551961
Rsp35_59 sp35_59 sp36_59 11.551961
Rsn35_59 sn35_59 sn36_59 11.551961
Rsp35_60 sp35_60 sp36_60 11.551961
Rsn35_60 sn35_60 sn36_60 11.551961
Rsp35_61 sp35_61 sp36_61 11.551961
Rsn35_61 sn35_61 sn36_61 11.551961
Rsp35_62 sp35_62 sp36_62 11.551961
Rsn35_62 sn35_62 sn36_62 11.551961
Rsp35_63 sp35_63 sp36_63 11.551961
Rsn35_63 sn35_63 sn36_63 11.551961
Rsp35_64 sp35_64 sp36_64 11.551961
Rsn35_64 sn35_64 sn36_64 11.551961
Rsp35_65 sp35_65 sp36_65 11.551961
Rsn35_65 sn35_65 sn36_65 11.551961
Rsp35_66 sp35_66 sp36_66 11.551961
Rsn35_66 sn35_66 sn36_66 11.551961
Rsp35_67 sp35_67 sp36_67 11.551961
Rsn35_67 sn35_67 sn36_67 11.551961
Rsp35_68 sp35_68 sp36_68 11.551961
Rsn35_68 sn35_68 sn36_68 11.551961
Rsp35_69 sp35_69 sp36_69 11.551961
Rsn35_69 sn35_69 sn36_69 11.551961
Rsp35_70 sp35_70 sp36_70 11.551961
Rsn35_70 sn35_70 sn36_70 11.551961
Rsp35_71 sp35_71 sp36_71 11.551961
Rsn35_71 sn35_71 sn36_71 11.551961
Rsp35_72 sp35_72 sp36_72 11.551961
Rsn35_72 sn35_72 sn36_72 11.551961
Rsp35_73 sp35_73 sp36_73 11.551961
Rsn35_73 sn35_73 sn36_73 11.551961
Rsp35_74 sp35_74 sp36_74 11.551961
Rsn35_74 sn35_74 sn36_74 11.551961
Rsp35_75 sp35_75 sp36_75 11.551961
Rsn35_75 sn35_75 sn36_75 11.551961
Rsp35_76 sp35_76 sp36_76 11.551961
Rsn35_76 sn35_76 sn36_76 11.551961
Rsp35_77 sp35_77 sp36_77 11.551961
Rsn35_77 sn35_77 sn36_77 11.551961
Rsp35_78 sp35_78 sp36_78 11.551961
Rsn35_78 sn35_78 sn36_78 11.551961
Rsp35_79 sp35_79 sp36_79 11.551961
Rsn35_79 sn35_79 sn36_79 11.551961
Rsp35_80 sp35_80 sp36_80 11.551961
Rsn35_80 sn35_80 sn36_80 11.551961
Rsp35_81 sp35_81 sp36_81 11.551961
Rsn35_81 sn35_81 sn36_81 11.551961
Rsp35_82 sp35_82 sp36_82 11.551961
Rsn35_82 sn35_82 sn36_82 11.551961
Rsp35_83 sp35_83 sp36_83 11.551961
Rsn35_83 sn35_83 sn36_83 11.551961
Rsp35_84 sp35_84 sp36_84 11.551961
Rsn35_84 sn35_84 sn36_84 11.551961
Rsp36_1 sp36_1 sp37_1 11.551961
Rsn36_1 sn36_1 sn37_1 11.551961
Rsp36_2 sp36_2 sp37_2 11.551961
Rsn36_2 sn36_2 sn37_2 11.551961
Rsp36_3 sp36_3 sp37_3 11.551961
Rsn36_3 sn36_3 sn37_3 11.551961
Rsp36_4 sp36_4 sp37_4 11.551961
Rsn36_4 sn36_4 sn37_4 11.551961
Rsp36_5 sp36_5 sp37_5 11.551961
Rsn36_5 sn36_5 sn37_5 11.551961
Rsp36_6 sp36_6 sp37_6 11.551961
Rsn36_6 sn36_6 sn37_6 11.551961
Rsp36_7 sp36_7 sp37_7 11.551961
Rsn36_7 sn36_7 sn37_7 11.551961
Rsp36_8 sp36_8 sp37_8 11.551961
Rsn36_8 sn36_8 sn37_8 11.551961
Rsp36_9 sp36_9 sp37_9 11.551961
Rsn36_9 sn36_9 sn37_9 11.551961
Rsp36_10 sp36_10 sp37_10 11.551961
Rsn36_10 sn36_10 sn37_10 11.551961
Rsp36_11 sp36_11 sp37_11 11.551961
Rsn36_11 sn36_11 sn37_11 11.551961
Rsp36_12 sp36_12 sp37_12 11.551961
Rsn36_12 sn36_12 sn37_12 11.551961
Rsp36_13 sp36_13 sp37_13 11.551961
Rsn36_13 sn36_13 sn37_13 11.551961
Rsp36_14 sp36_14 sp37_14 11.551961
Rsn36_14 sn36_14 sn37_14 11.551961
Rsp36_15 sp36_15 sp37_15 11.551961
Rsn36_15 sn36_15 sn37_15 11.551961
Rsp36_16 sp36_16 sp37_16 11.551961
Rsn36_16 sn36_16 sn37_16 11.551961
Rsp36_17 sp36_17 sp37_17 11.551961
Rsn36_17 sn36_17 sn37_17 11.551961
Rsp36_18 sp36_18 sp37_18 11.551961
Rsn36_18 sn36_18 sn37_18 11.551961
Rsp36_19 sp36_19 sp37_19 11.551961
Rsn36_19 sn36_19 sn37_19 11.551961
Rsp36_20 sp36_20 sp37_20 11.551961
Rsn36_20 sn36_20 sn37_20 11.551961
Rsp36_21 sp36_21 sp37_21 11.551961
Rsn36_21 sn36_21 sn37_21 11.551961
Rsp36_22 sp36_22 sp37_22 11.551961
Rsn36_22 sn36_22 sn37_22 11.551961
Rsp36_23 sp36_23 sp37_23 11.551961
Rsn36_23 sn36_23 sn37_23 11.551961
Rsp36_24 sp36_24 sp37_24 11.551961
Rsn36_24 sn36_24 sn37_24 11.551961
Rsp36_25 sp36_25 sp37_25 11.551961
Rsn36_25 sn36_25 sn37_25 11.551961
Rsp36_26 sp36_26 sp37_26 11.551961
Rsn36_26 sn36_26 sn37_26 11.551961
Rsp36_27 sp36_27 sp37_27 11.551961
Rsn36_27 sn36_27 sn37_27 11.551961
Rsp36_28 sp36_28 sp37_28 11.551961
Rsn36_28 sn36_28 sn37_28 11.551961
Rsp36_29 sp36_29 sp37_29 11.551961
Rsn36_29 sn36_29 sn37_29 11.551961
Rsp36_30 sp36_30 sp37_30 11.551961
Rsn36_30 sn36_30 sn37_30 11.551961
Rsp36_31 sp36_31 sp37_31 11.551961
Rsn36_31 sn36_31 sn37_31 11.551961
Rsp36_32 sp36_32 sp37_32 11.551961
Rsn36_32 sn36_32 sn37_32 11.551961
Rsp36_33 sp36_33 sp37_33 11.551961
Rsn36_33 sn36_33 sn37_33 11.551961
Rsp36_34 sp36_34 sp37_34 11.551961
Rsn36_34 sn36_34 sn37_34 11.551961
Rsp36_35 sp36_35 sp37_35 11.551961
Rsn36_35 sn36_35 sn37_35 11.551961
Rsp36_36 sp36_36 sp37_36 11.551961
Rsn36_36 sn36_36 sn37_36 11.551961
Rsp36_37 sp36_37 sp37_37 11.551961
Rsn36_37 sn36_37 sn37_37 11.551961
Rsp36_38 sp36_38 sp37_38 11.551961
Rsn36_38 sn36_38 sn37_38 11.551961
Rsp36_39 sp36_39 sp37_39 11.551961
Rsn36_39 sn36_39 sn37_39 11.551961
Rsp36_40 sp36_40 sp37_40 11.551961
Rsn36_40 sn36_40 sn37_40 11.551961
Rsp36_41 sp36_41 sp37_41 11.551961
Rsn36_41 sn36_41 sn37_41 11.551961
Rsp36_42 sp36_42 sp37_42 11.551961
Rsn36_42 sn36_42 sn37_42 11.551961
Rsp36_43 sp36_43 sp37_43 11.551961
Rsn36_43 sn36_43 sn37_43 11.551961
Rsp36_44 sp36_44 sp37_44 11.551961
Rsn36_44 sn36_44 sn37_44 11.551961
Rsp36_45 sp36_45 sp37_45 11.551961
Rsn36_45 sn36_45 sn37_45 11.551961
Rsp36_46 sp36_46 sp37_46 11.551961
Rsn36_46 sn36_46 sn37_46 11.551961
Rsp36_47 sp36_47 sp37_47 11.551961
Rsn36_47 sn36_47 sn37_47 11.551961
Rsp36_48 sp36_48 sp37_48 11.551961
Rsn36_48 sn36_48 sn37_48 11.551961
Rsp36_49 sp36_49 sp37_49 11.551961
Rsn36_49 sn36_49 sn37_49 11.551961
Rsp36_50 sp36_50 sp37_50 11.551961
Rsn36_50 sn36_50 sn37_50 11.551961
Rsp36_51 sp36_51 sp37_51 11.551961
Rsn36_51 sn36_51 sn37_51 11.551961
Rsp36_52 sp36_52 sp37_52 11.551961
Rsn36_52 sn36_52 sn37_52 11.551961
Rsp36_53 sp36_53 sp37_53 11.551961
Rsn36_53 sn36_53 sn37_53 11.551961
Rsp36_54 sp36_54 sp37_54 11.551961
Rsn36_54 sn36_54 sn37_54 11.551961
Rsp36_55 sp36_55 sp37_55 11.551961
Rsn36_55 sn36_55 sn37_55 11.551961
Rsp36_56 sp36_56 sp37_56 11.551961
Rsn36_56 sn36_56 sn37_56 11.551961
Rsp36_57 sp36_57 sp37_57 11.551961
Rsn36_57 sn36_57 sn37_57 11.551961
Rsp36_58 sp36_58 sp37_58 11.551961
Rsn36_58 sn36_58 sn37_58 11.551961
Rsp36_59 sp36_59 sp37_59 11.551961
Rsn36_59 sn36_59 sn37_59 11.551961
Rsp36_60 sp36_60 sp37_60 11.551961
Rsn36_60 sn36_60 sn37_60 11.551961
Rsp36_61 sp36_61 sp37_61 11.551961
Rsn36_61 sn36_61 sn37_61 11.551961
Rsp36_62 sp36_62 sp37_62 11.551961
Rsn36_62 sn36_62 sn37_62 11.551961
Rsp36_63 sp36_63 sp37_63 11.551961
Rsn36_63 sn36_63 sn37_63 11.551961
Rsp36_64 sp36_64 sp37_64 11.551961
Rsn36_64 sn36_64 sn37_64 11.551961
Rsp36_65 sp36_65 sp37_65 11.551961
Rsn36_65 sn36_65 sn37_65 11.551961
Rsp36_66 sp36_66 sp37_66 11.551961
Rsn36_66 sn36_66 sn37_66 11.551961
Rsp36_67 sp36_67 sp37_67 11.551961
Rsn36_67 sn36_67 sn37_67 11.551961
Rsp36_68 sp36_68 sp37_68 11.551961
Rsn36_68 sn36_68 sn37_68 11.551961
Rsp36_69 sp36_69 sp37_69 11.551961
Rsn36_69 sn36_69 sn37_69 11.551961
Rsp36_70 sp36_70 sp37_70 11.551961
Rsn36_70 sn36_70 sn37_70 11.551961
Rsp36_71 sp36_71 sp37_71 11.551961
Rsn36_71 sn36_71 sn37_71 11.551961
Rsp36_72 sp36_72 sp37_72 11.551961
Rsn36_72 sn36_72 sn37_72 11.551961
Rsp36_73 sp36_73 sp37_73 11.551961
Rsn36_73 sn36_73 sn37_73 11.551961
Rsp36_74 sp36_74 sp37_74 11.551961
Rsn36_74 sn36_74 sn37_74 11.551961
Rsp36_75 sp36_75 sp37_75 11.551961
Rsn36_75 sn36_75 sn37_75 11.551961
Rsp36_76 sp36_76 sp37_76 11.551961
Rsn36_76 sn36_76 sn37_76 11.551961
Rsp36_77 sp36_77 sp37_77 11.551961
Rsn36_77 sn36_77 sn37_77 11.551961
Rsp36_78 sp36_78 sp37_78 11.551961
Rsn36_78 sn36_78 sn37_78 11.551961
Rsp36_79 sp36_79 sp37_79 11.551961
Rsn36_79 sn36_79 sn37_79 11.551961
Rsp36_80 sp36_80 sp37_80 11.551961
Rsn36_80 sn36_80 sn37_80 11.551961
Rsp36_81 sp36_81 sp37_81 11.551961
Rsn36_81 sn36_81 sn37_81 11.551961
Rsp36_82 sp36_82 sp37_82 11.551961
Rsn36_82 sn36_82 sn37_82 11.551961
Rsp36_83 sp36_83 sp37_83 11.551961
Rsn36_83 sn36_83 sn37_83 11.551961
Rsp36_84 sp36_84 sp37_84 11.551961
Rsn36_84 sn36_84 sn37_84 11.551961
Rsp37_1 sp37_1 sp38_1 11.551961
Rsn37_1 sn37_1 sn38_1 11.551961
Rsp37_2 sp37_2 sp38_2 11.551961
Rsn37_2 sn37_2 sn38_2 11.551961
Rsp37_3 sp37_3 sp38_3 11.551961
Rsn37_3 sn37_3 sn38_3 11.551961
Rsp37_4 sp37_4 sp38_4 11.551961
Rsn37_4 sn37_4 sn38_4 11.551961
Rsp37_5 sp37_5 sp38_5 11.551961
Rsn37_5 sn37_5 sn38_5 11.551961
Rsp37_6 sp37_6 sp38_6 11.551961
Rsn37_6 sn37_6 sn38_6 11.551961
Rsp37_7 sp37_7 sp38_7 11.551961
Rsn37_7 sn37_7 sn38_7 11.551961
Rsp37_8 sp37_8 sp38_8 11.551961
Rsn37_8 sn37_8 sn38_8 11.551961
Rsp37_9 sp37_9 sp38_9 11.551961
Rsn37_9 sn37_9 sn38_9 11.551961
Rsp37_10 sp37_10 sp38_10 11.551961
Rsn37_10 sn37_10 sn38_10 11.551961
Rsp37_11 sp37_11 sp38_11 11.551961
Rsn37_11 sn37_11 sn38_11 11.551961
Rsp37_12 sp37_12 sp38_12 11.551961
Rsn37_12 sn37_12 sn38_12 11.551961
Rsp37_13 sp37_13 sp38_13 11.551961
Rsn37_13 sn37_13 sn38_13 11.551961
Rsp37_14 sp37_14 sp38_14 11.551961
Rsn37_14 sn37_14 sn38_14 11.551961
Rsp37_15 sp37_15 sp38_15 11.551961
Rsn37_15 sn37_15 sn38_15 11.551961
Rsp37_16 sp37_16 sp38_16 11.551961
Rsn37_16 sn37_16 sn38_16 11.551961
Rsp37_17 sp37_17 sp38_17 11.551961
Rsn37_17 sn37_17 sn38_17 11.551961
Rsp37_18 sp37_18 sp38_18 11.551961
Rsn37_18 sn37_18 sn38_18 11.551961
Rsp37_19 sp37_19 sp38_19 11.551961
Rsn37_19 sn37_19 sn38_19 11.551961
Rsp37_20 sp37_20 sp38_20 11.551961
Rsn37_20 sn37_20 sn38_20 11.551961
Rsp37_21 sp37_21 sp38_21 11.551961
Rsn37_21 sn37_21 sn38_21 11.551961
Rsp37_22 sp37_22 sp38_22 11.551961
Rsn37_22 sn37_22 sn38_22 11.551961
Rsp37_23 sp37_23 sp38_23 11.551961
Rsn37_23 sn37_23 sn38_23 11.551961
Rsp37_24 sp37_24 sp38_24 11.551961
Rsn37_24 sn37_24 sn38_24 11.551961
Rsp37_25 sp37_25 sp38_25 11.551961
Rsn37_25 sn37_25 sn38_25 11.551961
Rsp37_26 sp37_26 sp38_26 11.551961
Rsn37_26 sn37_26 sn38_26 11.551961
Rsp37_27 sp37_27 sp38_27 11.551961
Rsn37_27 sn37_27 sn38_27 11.551961
Rsp37_28 sp37_28 sp38_28 11.551961
Rsn37_28 sn37_28 sn38_28 11.551961
Rsp37_29 sp37_29 sp38_29 11.551961
Rsn37_29 sn37_29 sn38_29 11.551961
Rsp37_30 sp37_30 sp38_30 11.551961
Rsn37_30 sn37_30 sn38_30 11.551961
Rsp37_31 sp37_31 sp38_31 11.551961
Rsn37_31 sn37_31 sn38_31 11.551961
Rsp37_32 sp37_32 sp38_32 11.551961
Rsn37_32 sn37_32 sn38_32 11.551961
Rsp37_33 sp37_33 sp38_33 11.551961
Rsn37_33 sn37_33 sn38_33 11.551961
Rsp37_34 sp37_34 sp38_34 11.551961
Rsn37_34 sn37_34 sn38_34 11.551961
Rsp37_35 sp37_35 sp38_35 11.551961
Rsn37_35 sn37_35 sn38_35 11.551961
Rsp37_36 sp37_36 sp38_36 11.551961
Rsn37_36 sn37_36 sn38_36 11.551961
Rsp37_37 sp37_37 sp38_37 11.551961
Rsn37_37 sn37_37 sn38_37 11.551961
Rsp37_38 sp37_38 sp38_38 11.551961
Rsn37_38 sn37_38 sn38_38 11.551961
Rsp37_39 sp37_39 sp38_39 11.551961
Rsn37_39 sn37_39 sn38_39 11.551961
Rsp37_40 sp37_40 sp38_40 11.551961
Rsn37_40 sn37_40 sn38_40 11.551961
Rsp37_41 sp37_41 sp38_41 11.551961
Rsn37_41 sn37_41 sn38_41 11.551961
Rsp37_42 sp37_42 sp38_42 11.551961
Rsn37_42 sn37_42 sn38_42 11.551961
Rsp37_43 sp37_43 sp38_43 11.551961
Rsn37_43 sn37_43 sn38_43 11.551961
Rsp37_44 sp37_44 sp38_44 11.551961
Rsn37_44 sn37_44 sn38_44 11.551961
Rsp37_45 sp37_45 sp38_45 11.551961
Rsn37_45 sn37_45 sn38_45 11.551961
Rsp37_46 sp37_46 sp38_46 11.551961
Rsn37_46 sn37_46 sn38_46 11.551961
Rsp37_47 sp37_47 sp38_47 11.551961
Rsn37_47 sn37_47 sn38_47 11.551961
Rsp37_48 sp37_48 sp38_48 11.551961
Rsn37_48 sn37_48 sn38_48 11.551961
Rsp37_49 sp37_49 sp38_49 11.551961
Rsn37_49 sn37_49 sn38_49 11.551961
Rsp37_50 sp37_50 sp38_50 11.551961
Rsn37_50 sn37_50 sn38_50 11.551961
Rsp37_51 sp37_51 sp38_51 11.551961
Rsn37_51 sn37_51 sn38_51 11.551961
Rsp37_52 sp37_52 sp38_52 11.551961
Rsn37_52 sn37_52 sn38_52 11.551961
Rsp37_53 sp37_53 sp38_53 11.551961
Rsn37_53 sn37_53 sn38_53 11.551961
Rsp37_54 sp37_54 sp38_54 11.551961
Rsn37_54 sn37_54 sn38_54 11.551961
Rsp37_55 sp37_55 sp38_55 11.551961
Rsn37_55 sn37_55 sn38_55 11.551961
Rsp37_56 sp37_56 sp38_56 11.551961
Rsn37_56 sn37_56 sn38_56 11.551961
Rsp37_57 sp37_57 sp38_57 11.551961
Rsn37_57 sn37_57 sn38_57 11.551961
Rsp37_58 sp37_58 sp38_58 11.551961
Rsn37_58 sn37_58 sn38_58 11.551961
Rsp37_59 sp37_59 sp38_59 11.551961
Rsn37_59 sn37_59 sn38_59 11.551961
Rsp37_60 sp37_60 sp38_60 11.551961
Rsn37_60 sn37_60 sn38_60 11.551961
Rsp37_61 sp37_61 sp38_61 11.551961
Rsn37_61 sn37_61 sn38_61 11.551961
Rsp37_62 sp37_62 sp38_62 11.551961
Rsn37_62 sn37_62 sn38_62 11.551961
Rsp37_63 sp37_63 sp38_63 11.551961
Rsn37_63 sn37_63 sn38_63 11.551961
Rsp37_64 sp37_64 sp38_64 11.551961
Rsn37_64 sn37_64 sn38_64 11.551961
Rsp37_65 sp37_65 sp38_65 11.551961
Rsn37_65 sn37_65 sn38_65 11.551961
Rsp37_66 sp37_66 sp38_66 11.551961
Rsn37_66 sn37_66 sn38_66 11.551961
Rsp37_67 sp37_67 sp38_67 11.551961
Rsn37_67 sn37_67 sn38_67 11.551961
Rsp37_68 sp37_68 sp38_68 11.551961
Rsn37_68 sn37_68 sn38_68 11.551961
Rsp37_69 sp37_69 sp38_69 11.551961
Rsn37_69 sn37_69 sn38_69 11.551961
Rsp37_70 sp37_70 sp38_70 11.551961
Rsn37_70 sn37_70 sn38_70 11.551961
Rsp37_71 sp37_71 sp38_71 11.551961
Rsn37_71 sn37_71 sn38_71 11.551961
Rsp37_72 sp37_72 sp38_72 11.551961
Rsn37_72 sn37_72 sn38_72 11.551961
Rsp37_73 sp37_73 sp38_73 11.551961
Rsn37_73 sn37_73 sn38_73 11.551961
Rsp37_74 sp37_74 sp38_74 11.551961
Rsn37_74 sn37_74 sn38_74 11.551961
Rsp37_75 sp37_75 sp38_75 11.551961
Rsn37_75 sn37_75 sn38_75 11.551961
Rsp37_76 sp37_76 sp38_76 11.551961
Rsn37_76 sn37_76 sn38_76 11.551961
Rsp37_77 sp37_77 sp38_77 11.551961
Rsn37_77 sn37_77 sn38_77 11.551961
Rsp37_78 sp37_78 sp38_78 11.551961
Rsn37_78 sn37_78 sn38_78 11.551961
Rsp37_79 sp37_79 sp38_79 11.551961
Rsn37_79 sn37_79 sn38_79 11.551961
Rsp37_80 sp37_80 sp38_80 11.551961
Rsn37_80 sn37_80 sn38_80 11.551961
Rsp37_81 sp37_81 sp38_81 11.551961
Rsn37_81 sn37_81 sn38_81 11.551961
Rsp37_82 sp37_82 sp38_82 11.551961
Rsn37_82 sn37_82 sn38_82 11.551961
Rsp37_83 sp37_83 sp38_83 11.551961
Rsn37_83 sn37_83 sn38_83 11.551961
Rsp37_84 sp37_84 sp38_84 11.551961
Rsn37_84 sn37_84 sn38_84 11.551961
Rsp38_1 sp38_1 sp39_1 11.551961
Rsn38_1 sn38_1 sn39_1 11.551961
Rsp38_2 sp38_2 sp39_2 11.551961
Rsn38_2 sn38_2 sn39_2 11.551961
Rsp38_3 sp38_3 sp39_3 11.551961
Rsn38_3 sn38_3 sn39_3 11.551961
Rsp38_4 sp38_4 sp39_4 11.551961
Rsn38_4 sn38_4 sn39_4 11.551961
Rsp38_5 sp38_5 sp39_5 11.551961
Rsn38_5 sn38_5 sn39_5 11.551961
Rsp38_6 sp38_6 sp39_6 11.551961
Rsn38_6 sn38_6 sn39_6 11.551961
Rsp38_7 sp38_7 sp39_7 11.551961
Rsn38_7 sn38_7 sn39_7 11.551961
Rsp38_8 sp38_8 sp39_8 11.551961
Rsn38_8 sn38_8 sn39_8 11.551961
Rsp38_9 sp38_9 sp39_9 11.551961
Rsn38_9 sn38_9 sn39_9 11.551961
Rsp38_10 sp38_10 sp39_10 11.551961
Rsn38_10 sn38_10 sn39_10 11.551961
Rsp38_11 sp38_11 sp39_11 11.551961
Rsn38_11 sn38_11 sn39_11 11.551961
Rsp38_12 sp38_12 sp39_12 11.551961
Rsn38_12 sn38_12 sn39_12 11.551961
Rsp38_13 sp38_13 sp39_13 11.551961
Rsn38_13 sn38_13 sn39_13 11.551961
Rsp38_14 sp38_14 sp39_14 11.551961
Rsn38_14 sn38_14 sn39_14 11.551961
Rsp38_15 sp38_15 sp39_15 11.551961
Rsn38_15 sn38_15 sn39_15 11.551961
Rsp38_16 sp38_16 sp39_16 11.551961
Rsn38_16 sn38_16 sn39_16 11.551961
Rsp38_17 sp38_17 sp39_17 11.551961
Rsn38_17 sn38_17 sn39_17 11.551961
Rsp38_18 sp38_18 sp39_18 11.551961
Rsn38_18 sn38_18 sn39_18 11.551961
Rsp38_19 sp38_19 sp39_19 11.551961
Rsn38_19 sn38_19 sn39_19 11.551961
Rsp38_20 sp38_20 sp39_20 11.551961
Rsn38_20 sn38_20 sn39_20 11.551961
Rsp38_21 sp38_21 sp39_21 11.551961
Rsn38_21 sn38_21 sn39_21 11.551961
Rsp38_22 sp38_22 sp39_22 11.551961
Rsn38_22 sn38_22 sn39_22 11.551961
Rsp38_23 sp38_23 sp39_23 11.551961
Rsn38_23 sn38_23 sn39_23 11.551961
Rsp38_24 sp38_24 sp39_24 11.551961
Rsn38_24 sn38_24 sn39_24 11.551961
Rsp38_25 sp38_25 sp39_25 11.551961
Rsn38_25 sn38_25 sn39_25 11.551961
Rsp38_26 sp38_26 sp39_26 11.551961
Rsn38_26 sn38_26 sn39_26 11.551961
Rsp38_27 sp38_27 sp39_27 11.551961
Rsn38_27 sn38_27 sn39_27 11.551961
Rsp38_28 sp38_28 sp39_28 11.551961
Rsn38_28 sn38_28 sn39_28 11.551961
Rsp38_29 sp38_29 sp39_29 11.551961
Rsn38_29 sn38_29 sn39_29 11.551961
Rsp38_30 sp38_30 sp39_30 11.551961
Rsn38_30 sn38_30 sn39_30 11.551961
Rsp38_31 sp38_31 sp39_31 11.551961
Rsn38_31 sn38_31 sn39_31 11.551961
Rsp38_32 sp38_32 sp39_32 11.551961
Rsn38_32 sn38_32 sn39_32 11.551961
Rsp38_33 sp38_33 sp39_33 11.551961
Rsn38_33 sn38_33 sn39_33 11.551961
Rsp38_34 sp38_34 sp39_34 11.551961
Rsn38_34 sn38_34 sn39_34 11.551961
Rsp38_35 sp38_35 sp39_35 11.551961
Rsn38_35 sn38_35 sn39_35 11.551961
Rsp38_36 sp38_36 sp39_36 11.551961
Rsn38_36 sn38_36 sn39_36 11.551961
Rsp38_37 sp38_37 sp39_37 11.551961
Rsn38_37 sn38_37 sn39_37 11.551961
Rsp38_38 sp38_38 sp39_38 11.551961
Rsn38_38 sn38_38 sn39_38 11.551961
Rsp38_39 sp38_39 sp39_39 11.551961
Rsn38_39 sn38_39 sn39_39 11.551961
Rsp38_40 sp38_40 sp39_40 11.551961
Rsn38_40 sn38_40 sn39_40 11.551961
Rsp38_41 sp38_41 sp39_41 11.551961
Rsn38_41 sn38_41 sn39_41 11.551961
Rsp38_42 sp38_42 sp39_42 11.551961
Rsn38_42 sn38_42 sn39_42 11.551961
Rsp38_43 sp38_43 sp39_43 11.551961
Rsn38_43 sn38_43 sn39_43 11.551961
Rsp38_44 sp38_44 sp39_44 11.551961
Rsn38_44 sn38_44 sn39_44 11.551961
Rsp38_45 sp38_45 sp39_45 11.551961
Rsn38_45 sn38_45 sn39_45 11.551961
Rsp38_46 sp38_46 sp39_46 11.551961
Rsn38_46 sn38_46 sn39_46 11.551961
Rsp38_47 sp38_47 sp39_47 11.551961
Rsn38_47 sn38_47 sn39_47 11.551961
Rsp38_48 sp38_48 sp39_48 11.551961
Rsn38_48 sn38_48 sn39_48 11.551961
Rsp38_49 sp38_49 sp39_49 11.551961
Rsn38_49 sn38_49 sn39_49 11.551961
Rsp38_50 sp38_50 sp39_50 11.551961
Rsn38_50 sn38_50 sn39_50 11.551961
Rsp38_51 sp38_51 sp39_51 11.551961
Rsn38_51 sn38_51 sn39_51 11.551961
Rsp38_52 sp38_52 sp39_52 11.551961
Rsn38_52 sn38_52 sn39_52 11.551961
Rsp38_53 sp38_53 sp39_53 11.551961
Rsn38_53 sn38_53 sn39_53 11.551961
Rsp38_54 sp38_54 sp39_54 11.551961
Rsn38_54 sn38_54 sn39_54 11.551961
Rsp38_55 sp38_55 sp39_55 11.551961
Rsn38_55 sn38_55 sn39_55 11.551961
Rsp38_56 sp38_56 sp39_56 11.551961
Rsn38_56 sn38_56 sn39_56 11.551961
Rsp38_57 sp38_57 sp39_57 11.551961
Rsn38_57 sn38_57 sn39_57 11.551961
Rsp38_58 sp38_58 sp39_58 11.551961
Rsn38_58 sn38_58 sn39_58 11.551961
Rsp38_59 sp38_59 sp39_59 11.551961
Rsn38_59 sn38_59 sn39_59 11.551961
Rsp38_60 sp38_60 sp39_60 11.551961
Rsn38_60 sn38_60 sn39_60 11.551961
Rsp38_61 sp38_61 sp39_61 11.551961
Rsn38_61 sn38_61 sn39_61 11.551961
Rsp38_62 sp38_62 sp39_62 11.551961
Rsn38_62 sn38_62 sn39_62 11.551961
Rsp38_63 sp38_63 sp39_63 11.551961
Rsn38_63 sn38_63 sn39_63 11.551961
Rsp38_64 sp38_64 sp39_64 11.551961
Rsn38_64 sn38_64 sn39_64 11.551961
Rsp38_65 sp38_65 sp39_65 11.551961
Rsn38_65 sn38_65 sn39_65 11.551961
Rsp38_66 sp38_66 sp39_66 11.551961
Rsn38_66 sn38_66 sn39_66 11.551961
Rsp38_67 sp38_67 sp39_67 11.551961
Rsn38_67 sn38_67 sn39_67 11.551961
Rsp38_68 sp38_68 sp39_68 11.551961
Rsn38_68 sn38_68 sn39_68 11.551961
Rsp38_69 sp38_69 sp39_69 11.551961
Rsn38_69 sn38_69 sn39_69 11.551961
Rsp38_70 sp38_70 sp39_70 11.551961
Rsn38_70 sn38_70 sn39_70 11.551961
Rsp38_71 sp38_71 sp39_71 11.551961
Rsn38_71 sn38_71 sn39_71 11.551961
Rsp38_72 sp38_72 sp39_72 11.551961
Rsn38_72 sn38_72 sn39_72 11.551961
Rsp38_73 sp38_73 sp39_73 11.551961
Rsn38_73 sn38_73 sn39_73 11.551961
Rsp38_74 sp38_74 sp39_74 11.551961
Rsn38_74 sn38_74 sn39_74 11.551961
Rsp38_75 sp38_75 sp39_75 11.551961
Rsn38_75 sn38_75 sn39_75 11.551961
Rsp38_76 sp38_76 sp39_76 11.551961
Rsn38_76 sn38_76 sn39_76 11.551961
Rsp38_77 sp38_77 sp39_77 11.551961
Rsn38_77 sn38_77 sn39_77 11.551961
Rsp38_78 sp38_78 sp39_78 11.551961
Rsn38_78 sn38_78 sn39_78 11.551961
Rsp38_79 sp38_79 sp39_79 11.551961
Rsn38_79 sn38_79 sn39_79 11.551961
Rsp38_80 sp38_80 sp39_80 11.551961
Rsn38_80 sn38_80 sn39_80 11.551961
Rsp38_81 sp38_81 sp39_81 11.551961
Rsn38_81 sn38_81 sn39_81 11.551961
Rsp38_82 sp38_82 sp39_82 11.551961
Rsn38_82 sn38_82 sn39_82 11.551961
Rsp38_83 sp38_83 sp39_83 11.551961
Rsn38_83 sn38_83 sn39_83 11.551961
Rsp38_84 sp38_84 sp39_84 11.551961
Rsn38_84 sn38_84 sn39_84 11.551961
Rsp39_1 sp39_1 sp40_1 11.551961
Rsn39_1 sn39_1 sn40_1 11.551961
Rsp39_2 sp39_2 sp40_2 11.551961
Rsn39_2 sn39_2 sn40_2 11.551961
Rsp39_3 sp39_3 sp40_3 11.551961
Rsn39_3 sn39_3 sn40_3 11.551961
Rsp39_4 sp39_4 sp40_4 11.551961
Rsn39_4 sn39_4 sn40_4 11.551961
Rsp39_5 sp39_5 sp40_5 11.551961
Rsn39_5 sn39_5 sn40_5 11.551961
Rsp39_6 sp39_6 sp40_6 11.551961
Rsn39_6 sn39_6 sn40_6 11.551961
Rsp39_7 sp39_7 sp40_7 11.551961
Rsn39_7 sn39_7 sn40_7 11.551961
Rsp39_8 sp39_8 sp40_8 11.551961
Rsn39_8 sn39_8 sn40_8 11.551961
Rsp39_9 sp39_9 sp40_9 11.551961
Rsn39_9 sn39_9 sn40_9 11.551961
Rsp39_10 sp39_10 sp40_10 11.551961
Rsn39_10 sn39_10 sn40_10 11.551961
Rsp39_11 sp39_11 sp40_11 11.551961
Rsn39_11 sn39_11 sn40_11 11.551961
Rsp39_12 sp39_12 sp40_12 11.551961
Rsn39_12 sn39_12 sn40_12 11.551961
Rsp39_13 sp39_13 sp40_13 11.551961
Rsn39_13 sn39_13 sn40_13 11.551961
Rsp39_14 sp39_14 sp40_14 11.551961
Rsn39_14 sn39_14 sn40_14 11.551961
Rsp39_15 sp39_15 sp40_15 11.551961
Rsn39_15 sn39_15 sn40_15 11.551961
Rsp39_16 sp39_16 sp40_16 11.551961
Rsn39_16 sn39_16 sn40_16 11.551961
Rsp39_17 sp39_17 sp40_17 11.551961
Rsn39_17 sn39_17 sn40_17 11.551961
Rsp39_18 sp39_18 sp40_18 11.551961
Rsn39_18 sn39_18 sn40_18 11.551961
Rsp39_19 sp39_19 sp40_19 11.551961
Rsn39_19 sn39_19 sn40_19 11.551961
Rsp39_20 sp39_20 sp40_20 11.551961
Rsn39_20 sn39_20 sn40_20 11.551961
Rsp39_21 sp39_21 sp40_21 11.551961
Rsn39_21 sn39_21 sn40_21 11.551961
Rsp39_22 sp39_22 sp40_22 11.551961
Rsn39_22 sn39_22 sn40_22 11.551961
Rsp39_23 sp39_23 sp40_23 11.551961
Rsn39_23 sn39_23 sn40_23 11.551961
Rsp39_24 sp39_24 sp40_24 11.551961
Rsn39_24 sn39_24 sn40_24 11.551961
Rsp39_25 sp39_25 sp40_25 11.551961
Rsn39_25 sn39_25 sn40_25 11.551961
Rsp39_26 sp39_26 sp40_26 11.551961
Rsn39_26 sn39_26 sn40_26 11.551961
Rsp39_27 sp39_27 sp40_27 11.551961
Rsn39_27 sn39_27 sn40_27 11.551961
Rsp39_28 sp39_28 sp40_28 11.551961
Rsn39_28 sn39_28 sn40_28 11.551961
Rsp39_29 sp39_29 sp40_29 11.551961
Rsn39_29 sn39_29 sn40_29 11.551961
Rsp39_30 sp39_30 sp40_30 11.551961
Rsn39_30 sn39_30 sn40_30 11.551961
Rsp39_31 sp39_31 sp40_31 11.551961
Rsn39_31 sn39_31 sn40_31 11.551961
Rsp39_32 sp39_32 sp40_32 11.551961
Rsn39_32 sn39_32 sn40_32 11.551961
Rsp39_33 sp39_33 sp40_33 11.551961
Rsn39_33 sn39_33 sn40_33 11.551961
Rsp39_34 sp39_34 sp40_34 11.551961
Rsn39_34 sn39_34 sn40_34 11.551961
Rsp39_35 sp39_35 sp40_35 11.551961
Rsn39_35 sn39_35 sn40_35 11.551961
Rsp39_36 sp39_36 sp40_36 11.551961
Rsn39_36 sn39_36 sn40_36 11.551961
Rsp39_37 sp39_37 sp40_37 11.551961
Rsn39_37 sn39_37 sn40_37 11.551961
Rsp39_38 sp39_38 sp40_38 11.551961
Rsn39_38 sn39_38 sn40_38 11.551961
Rsp39_39 sp39_39 sp40_39 11.551961
Rsn39_39 sn39_39 sn40_39 11.551961
Rsp39_40 sp39_40 sp40_40 11.551961
Rsn39_40 sn39_40 sn40_40 11.551961
Rsp39_41 sp39_41 sp40_41 11.551961
Rsn39_41 sn39_41 sn40_41 11.551961
Rsp39_42 sp39_42 sp40_42 11.551961
Rsn39_42 sn39_42 sn40_42 11.551961
Rsp39_43 sp39_43 sp40_43 11.551961
Rsn39_43 sn39_43 sn40_43 11.551961
Rsp39_44 sp39_44 sp40_44 11.551961
Rsn39_44 sn39_44 sn40_44 11.551961
Rsp39_45 sp39_45 sp40_45 11.551961
Rsn39_45 sn39_45 sn40_45 11.551961
Rsp39_46 sp39_46 sp40_46 11.551961
Rsn39_46 sn39_46 sn40_46 11.551961
Rsp39_47 sp39_47 sp40_47 11.551961
Rsn39_47 sn39_47 sn40_47 11.551961
Rsp39_48 sp39_48 sp40_48 11.551961
Rsn39_48 sn39_48 sn40_48 11.551961
Rsp39_49 sp39_49 sp40_49 11.551961
Rsn39_49 sn39_49 sn40_49 11.551961
Rsp39_50 sp39_50 sp40_50 11.551961
Rsn39_50 sn39_50 sn40_50 11.551961
Rsp39_51 sp39_51 sp40_51 11.551961
Rsn39_51 sn39_51 sn40_51 11.551961
Rsp39_52 sp39_52 sp40_52 11.551961
Rsn39_52 sn39_52 sn40_52 11.551961
Rsp39_53 sp39_53 sp40_53 11.551961
Rsn39_53 sn39_53 sn40_53 11.551961
Rsp39_54 sp39_54 sp40_54 11.551961
Rsn39_54 sn39_54 sn40_54 11.551961
Rsp39_55 sp39_55 sp40_55 11.551961
Rsn39_55 sn39_55 sn40_55 11.551961
Rsp39_56 sp39_56 sp40_56 11.551961
Rsn39_56 sn39_56 sn40_56 11.551961
Rsp39_57 sp39_57 sp40_57 11.551961
Rsn39_57 sn39_57 sn40_57 11.551961
Rsp39_58 sp39_58 sp40_58 11.551961
Rsn39_58 sn39_58 sn40_58 11.551961
Rsp39_59 sp39_59 sp40_59 11.551961
Rsn39_59 sn39_59 sn40_59 11.551961
Rsp39_60 sp39_60 sp40_60 11.551961
Rsn39_60 sn39_60 sn40_60 11.551961
Rsp39_61 sp39_61 sp40_61 11.551961
Rsn39_61 sn39_61 sn40_61 11.551961
Rsp39_62 sp39_62 sp40_62 11.551961
Rsn39_62 sn39_62 sn40_62 11.551961
Rsp39_63 sp39_63 sp40_63 11.551961
Rsn39_63 sn39_63 sn40_63 11.551961
Rsp39_64 sp39_64 sp40_64 11.551961
Rsn39_64 sn39_64 sn40_64 11.551961
Rsp39_65 sp39_65 sp40_65 11.551961
Rsn39_65 sn39_65 sn40_65 11.551961
Rsp39_66 sp39_66 sp40_66 11.551961
Rsn39_66 sn39_66 sn40_66 11.551961
Rsp39_67 sp39_67 sp40_67 11.551961
Rsn39_67 sn39_67 sn40_67 11.551961
Rsp39_68 sp39_68 sp40_68 11.551961
Rsn39_68 sn39_68 sn40_68 11.551961
Rsp39_69 sp39_69 sp40_69 11.551961
Rsn39_69 sn39_69 sn40_69 11.551961
Rsp39_70 sp39_70 sp40_70 11.551961
Rsn39_70 sn39_70 sn40_70 11.551961
Rsp39_71 sp39_71 sp40_71 11.551961
Rsn39_71 sn39_71 sn40_71 11.551961
Rsp39_72 sp39_72 sp40_72 11.551961
Rsn39_72 sn39_72 sn40_72 11.551961
Rsp39_73 sp39_73 sp40_73 11.551961
Rsn39_73 sn39_73 sn40_73 11.551961
Rsp39_74 sp39_74 sp40_74 11.551961
Rsn39_74 sn39_74 sn40_74 11.551961
Rsp39_75 sp39_75 sp40_75 11.551961
Rsn39_75 sn39_75 sn40_75 11.551961
Rsp39_76 sp39_76 sp40_76 11.551961
Rsn39_76 sn39_76 sn40_76 11.551961
Rsp39_77 sp39_77 sp40_77 11.551961
Rsn39_77 sn39_77 sn40_77 11.551961
Rsp39_78 sp39_78 sp40_78 11.551961
Rsn39_78 sn39_78 sn40_78 11.551961
Rsp39_79 sp39_79 sp40_79 11.551961
Rsn39_79 sn39_79 sn40_79 11.551961
Rsp39_80 sp39_80 sp40_80 11.551961
Rsn39_80 sn39_80 sn40_80 11.551961
Rsp39_81 sp39_81 sp40_81 11.551961
Rsn39_81 sn39_81 sn40_81 11.551961
Rsp39_82 sp39_82 sp40_82 11.551961
Rsn39_82 sn39_82 sn40_82 11.551961
Rsp39_83 sp39_83 sp40_83 11.551961
Rsn39_83 sn39_83 sn40_83 11.551961
Rsp39_84 sp39_84 sp40_84 11.551961
Rsn39_84 sn39_84 sn40_84 11.551961
Rsp40_1 sp40_1 sp41_1 11.551961
Rsn40_1 sn40_1 sn41_1 11.551961
Rsp40_2 sp40_2 sp41_2 11.551961
Rsn40_2 sn40_2 sn41_2 11.551961
Rsp40_3 sp40_3 sp41_3 11.551961
Rsn40_3 sn40_3 sn41_3 11.551961
Rsp40_4 sp40_4 sp41_4 11.551961
Rsn40_4 sn40_4 sn41_4 11.551961
Rsp40_5 sp40_5 sp41_5 11.551961
Rsn40_5 sn40_5 sn41_5 11.551961
Rsp40_6 sp40_6 sp41_6 11.551961
Rsn40_6 sn40_6 sn41_6 11.551961
Rsp40_7 sp40_7 sp41_7 11.551961
Rsn40_7 sn40_7 sn41_7 11.551961
Rsp40_8 sp40_8 sp41_8 11.551961
Rsn40_8 sn40_8 sn41_8 11.551961
Rsp40_9 sp40_9 sp41_9 11.551961
Rsn40_9 sn40_9 sn41_9 11.551961
Rsp40_10 sp40_10 sp41_10 11.551961
Rsn40_10 sn40_10 sn41_10 11.551961
Rsp40_11 sp40_11 sp41_11 11.551961
Rsn40_11 sn40_11 sn41_11 11.551961
Rsp40_12 sp40_12 sp41_12 11.551961
Rsn40_12 sn40_12 sn41_12 11.551961
Rsp40_13 sp40_13 sp41_13 11.551961
Rsn40_13 sn40_13 sn41_13 11.551961
Rsp40_14 sp40_14 sp41_14 11.551961
Rsn40_14 sn40_14 sn41_14 11.551961
Rsp40_15 sp40_15 sp41_15 11.551961
Rsn40_15 sn40_15 sn41_15 11.551961
Rsp40_16 sp40_16 sp41_16 11.551961
Rsn40_16 sn40_16 sn41_16 11.551961
Rsp40_17 sp40_17 sp41_17 11.551961
Rsn40_17 sn40_17 sn41_17 11.551961
Rsp40_18 sp40_18 sp41_18 11.551961
Rsn40_18 sn40_18 sn41_18 11.551961
Rsp40_19 sp40_19 sp41_19 11.551961
Rsn40_19 sn40_19 sn41_19 11.551961
Rsp40_20 sp40_20 sp41_20 11.551961
Rsn40_20 sn40_20 sn41_20 11.551961
Rsp40_21 sp40_21 sp41_21 11.551961
Rsn40_21 sn40_21 sn41_21 11.551961
Rsp40_22 sp40_22 sp41_22 11.551961
Rsn40_22 sn40_22 sn41_22 11.551961
Rsp40_23 sp40_23 sp41_23 11.551961
Rsn40_23 sn40_23 sn41_23 11.551961
Rsp40_24 sp40_24 sp41_24 11.551961
Rsn40_24 sn40_24 sn41_24 11.551961
Rsp40_25 sp40_25 sp41_25 11.551961
Rsn40_25 sn40_25 sn41_25 11.551961
Rsp40_26 sp40_26 sp41_26 11.551961
Rsn40_26 sn40_26 sn41_26 11.551961
Rsp40_27 sp40_27 sp41_27 11.551961
Rsn40_27 sn40_27 sn41_27 11.551961
Rsp40_28 sp40_28 sp41_28 11.551961
Rsn40_28 sn40_28 sn41_28 11.551961
Rsp40_29 sp40_29 sp41_29 11.551961
Rsn40_29 sn40_29 sn41_29 11.551961
Rsp40_30 sp40_30 sp41_30 11.551961
Rsn40_30 sn40_30 sn41_30 11.551961
Rsp40_31 sp40_31 sp41_31 11.551961
Rsn40_31 sn40_31 sn41_31 11.551961
Rsp40_32 sp40_32 sp41_32 11.551961
Rsn40_32 sn40_32 sn41_32 11.551961
Rsp40_33 sp40_33 sp41_33 11.551961
Rsn40_33 sn40_33 sn41_33 11.551961
Rsp40_34 sp40_34 sp41_34 11.551961
Rsn40_34 sn40_34 sn41_34 11.551961
Rsp40_35 sp40_35 sp41_35 11.551961
Rsn40_35 sn40_35 sn41_35 11.551961
Rsp40_36 sp40_36 sp41_36 11.551961
Rsn40_36 sn40_36 sn41_36 11.551961
Rsp40_37 sp40_37 sp41_37 11.551961
Rsn40_37 sn40_37 sn41_37 11.551961
Rsp40_38 sp40_38 sp41_38 11.551961
Rsn40_38 sn40_38 sn41_38 11.551961
Rsp40_39 sp40_39 sp41_39 11.551961
Rsn40_39 sn40_39 sn41_39 11.551961
Rsp40_40 sp40_40 sp41_40 11.551961
Rsn40_40 sn40_40 sn41_40 11.551961
Rsp40_41 sp40_41 sp41_41 11.551961
Rsn40_41 sn40_41 sn41_41 11.551961
Rsp40_42 sp40_42 sp41_42 11.551961
Rsn40_42 sn40_42 sn41_42 11.551961
Rsp40_43 sp40_43 sp41_43 11.551961
Rsn40_43 sn40_43 sn41_43 11.551961
Rsp40_44 sp40_44 sp41_44 11.551961
Rsn40_44 sn40_44 sn41_44 11.551961
Rsp40_45 sp40_45 sp41_45 11.551961
Rsn40_45 sn40_45 sn41_45 11.551961
Rsp40_46 sp40_46 sp41_46 11.551961
Rsn40_46 sn40_46 sn41_46 11.551961
Rsp40_47 sp40_47 sp41_47 11.551961
Rsn40_47 sn40_47 sn41_47 11.551961
Rsp40_48 sp40_48 sp41_48 11.551961
Rsn40_48 sn40_48 sn41_48 11.551961
Rsp40_49 sp40_49 sp41_49 11.551961
Rsn40_49 sn40_49 sn41_49 11.551961
Rsp40_50 sp40_50 sp41_50 11.551961
Rsn40_50 sn40_50 sn41_50 11.551961
Rsp40_51 sp40_51 sp41_51 11.551961
Rsn40_51 sn40_51 sn41_51 11.551961
Rsp40_52 sp40_52 sp41_52 11.551961
Rsn40_52 sn40_52 sn41_52 11.551961
Rsp40_53 sp40_53 sp41_53 11.551961
Rsn40_53 sn40_53 sn41_53 11.551961
Rsp40_54 sp40_54 sp41_54 11.551961
Rsn40_54 sn40_54 sn41_54 11.551961
Rsp40_55 sp40_55 sp41_55 11.551961
Rsn40_55 sn40_55 sn41_55 11.551961
Rsp40_56 sp40_56 sp41_56 11.551961
Rsn40_56 sn40_56 sn41_56 11.551961
Rsp40_57 sp40_57 sp41_57 11.551961
Rsn40_57 sn40_57 sn41_57 11.551961
Rsp40_58 sp40_58 sp41_58 11.551961
Rsn40_58 sn40_58 sn41_58 11.551961
Rsp40_59 sp40_59 sp41_59 11.551961
Rsn40_59 sn40_59 sn41_59 11.551961
Rsp40_60 sp40_60 sp41_60 11.551961
Rsn40_60 sn40_60 sn41_60 11.551961
Rsp40_61 sp40_61 sp41_61 11.551961
Rsn40_61 sn40_61 sn41_61 11.551961
Rsp40_62 sp40_62 sp41_62 11.551961
Rsn40_62 sn40_62 sn41_62 11.551961
Rsp40_63 sp40_63 sp41_63 11.551961
Rsn40_63 sn40_63 sn41_63 11.551961
Rsp40_64 sp40_64 sp41_64 11.551961
Rsn40_64 sn40_64 sn41_64 11.551961
Rsp40_65 sp40_65 sp41_65 11.551961
Rsn40_65 sn40_65 sn41_65 11.551961
Rsp40_66 sp40_66 sp41_66 11.551961
Rsn40_66 sn40_66 sn41_66 11.551961
Rsp40_67 sp40_67 sp41_67 11.551961
Rsn40_67 sn40_67 sn41_67 11.551961
Rsp40_68 sp40_68 sp41_68 11.551961
Rsn40_68 sn40_68 sn41_68 11.551961
Rsp40_69 sp40_69 sp41_69 11.551961
Rsn40_69 sn40_69 sn41_69 11.551961
Rsp40_70 sp40_70 sp41_70 11.551961
Rsn40_70 sn40_70 sn41_70 11.551961
Rsp40_71 sp40_71 sp41_71 11.551961
Rsn40_71 sn40_71 sn41_71 11.551961
Rsp40_72 sp40_72 sp41_72 11.551961
Rsn40_72 sn40_72 sn41_72 11.551961
Rsp40_73 sp40_73 sp41_73 11.551961
Rsn40_73 sn40_73 sn41_73 11.551961
Rsp40_74 sp40_74 sp41_74 11.551961
Rsn40_74 sn40_74 sn41_74 11.551961
Rsp40_75 sp40_75 sp41_75 11.551961
Rsn40_75 sn40_75 sn41_75 11.551961
Rsp40_76 sp40_76 sp41_76 11.551961
Rsn40_76 sn40_76 sn41_76 11.551961
Rsp40_77 sp40_77 sp41_77 11.551961
Rsn40_77 sn40_77 sn41_77 11.551961
Rsp40_78 sp40_78 sp41_78 11.551961
Rsn40_78 sn40_78 sn41_78 11.551961
Rsp40_79 sp40_79 sp41_79 11.551961
Rsn40_79 sn40_79 sn41_79 11.551961
Rsp40_80 sp40_80 sp41_80 11.551961
Rsn40_80 sn40_80 sn41_80 11.551961
Rsp40_81 sp40_81 sp41_81 11.551961
Rsn40_81 sn40_81 sn41_81 11.551961
Rsp40_82 sp40_82 sp41_82 11.551961
Rsn40_82 sn40_82 sn41_82 11.551961
Rsp40_83 sp40_83 sp41_83 11.551961
Rsn40_83 sn40_83 sn41_83 11.551961
Rsp40_84 sp40_84 sp41_84 11.551961
Rsn40_84 sn40_84 sn41_84 11.551961
Rsp41_1 sp41_1 sp42_1 11.551961
Rsn41_1 sn41_1 sn42_1 11.551961
Rsp41_2 sp41_2 sp42_2 11.551961
Rsn41_2 sn41_2 sn42_2 11.551961
Rsp41_3 sp41_3 sp42_3 11.551961
Rsn41_3 sn41_3 sn42_3 11.551961
Rsp41_4 sp41_4 sp42_4 11.551961
Rsn41_4 sn41_4 sn42_4 11.551961
Rsp41_5 sp41_5 sp42_5 11.551961
Rsn41_5 sn41_5 sn42_5 11.551961
Rsp41_6 sp41_6 sp42_6 11.551961
Rsn41_6 sn41_6 sn42_6 11.551961
Rsp41_7 sp41_7 sp42_7 11.551961
Rsn41_7 sn41_7 sn42_7 11.551961
Rsp41_8 sp41_8 sp42_8 11.551961
Rsn41_8 sn41_8 sn42_8 11.551961
Rsp41_9 sp41_9 sp42_9 11.551961
Rsn41_9 sn41_9 sn42_9 11.551961
Rsp41_10 sp41_10 sp42_10 11.551961
Rsn41_10 sn41_10 sn42_10 11.551961
Rsp41_11 sp41_11 sp42_11 11.551961
Rsn41_11 sn41_11 sn42_11 11.551961
Rsp41_12 sp41_12 sp42_12 11.551961
Rsn41_12 sn41_12 sn42_12 11.551961
Rsp41_13 sp41_13 sp42_13 11.551961
Rsn41_13 sn41_13 sn42_13 11.551961
Rsp41_14 sp41_14 sp42_14 11.551961
Rsn41_14 sn41_14 sn42_14 11.551961
Rsp41_15 sp41_15 sp42_15 11.551961
Rsn41_15 sn41_15 sn42_15 11.551961
Rsp41_16 sp41_16 sp42_16 11.551961
Rsn41_16 sn41_16 sn42_16 11.551961
Rsp41_17 sp41_17 sp42_17 11.551961
Rsn41_17 sn41_17 sn42_17 11.551961
Rsp41_18 sp41_18 sp42_18 11.551961
Rsn41_18 sn41_18 sn42_18 11.551961
Rsp41_19 sp41_19 sp42_19 11.551961
Rsn41_19 sn41_19 sn42_19 11.551961
Rsp41_20 sp41_20 sp42_20 11.551961
Rsn41_20 sn41_20 sn42_20 11.551961
Rsp41_21 sp41_21 sp42_21 11.551961
Rsn41_21 sn41_21 sn42_21 11.551961
Rsp41_22 sp41_22 sp42_22 11.551961
Rsn41_22 sn41_22 sn42_22 11.551961
Rsp41_23 sp41_23 sp42_23 11.551961
Rsn41_23 sn41_23 sn42_23 11.551961
Rsp41_24 sp41_24 sp42_24 11.551961
Rsn41_24 sn41_24 sn42_24 11.551961
Rsp41_25 sp41_25 sp42_25 11.551961
Rsn41_25 sn41_25 sn42_25 11.551961
Rsp41_26 sp41_26 sp42_26 11.551961
Rsn41_26 sn41_26 sn42_26 11.551961
Rsp41_27 sp41_27 sp42_27 11.551961
Rsn41_27 sn41_27 sn42_27 11.551961
Rsp41_28 sp41_28 sp42_28 11.551961
Rsn41_28 sn41_28 sn42_28 11.551961
Rsp41_29 sp41_29 sp42_29 11.551961
Rsn41_29 sn41_29 sn42_29 11.551961
Rsp41_30 sp41_30 sp42_30 11.551961
Rsn41_30 sn41_30 sn42_30 11.551961
Rsp41_31 sp41_31 sp42_31 11.551961
Rsn41_31 sn41_31 sn42_31 11.551961
Rsp41_32 sp41_32 sp42_32 11.551961
Rsn41_32 sn41_32 sn42_32 11.551961
Rsp41_33 sp41_33 sp42_33 11.551961
Rsn41_33 sn41_33 sn42_33 11.551961
Rsp41_34 sp41_34 sp42_34 11.551961
Rsn41_34 sn41_34 sn42_34 11.551961
Rsp41_35 sp41_35 sp42_35 11.551961
Rsn41_35 sn41_35 sn42_35 11.551961
Rsp41_36 sp41_36 sp42_36 11.551961
Rsn41_36 sn41_36 sn42_36 11.551961
Rsp41_37 sp41_37 sp42_37 11.551961
Rsn41_37 sn41_37 sn42_37 11.551961
Rsp41_38 sp41_38 sp42_38 11.551961
Rsn41_38 sn41_38 sn42_38 11.551961
Rsp41_39 sp41_39 sp42_39 11.551961
Rsn41_39 sn41_39 sn42_39 11.551961
Rsp41_40 sp41_40 sp42_40 11.551961
Rsn41_40 sn41_40 sn42_40 11.551961
Rsp41_41 sp41_41 sp42_41 11.551961
Rsn41_41 sn41_41 sn42_41 11.551961
Rsp41_42 sp41_42 sp42_42 11.551961
Rsn41_42 sn41_42 sn42_42 11.551961
Rsp41_43 sp41_43 sp42_43 11.551961
Rsn41_43 sn41_43 sn42_43 11.551961
Rsp41_44 sp41_44 sp42_44 11.551961
Rsn41_44 sn41_44 sn42_44 11.551961
Rsp41_45 sp41_45 sp42_45 11.551961
Rsn41_45 sn41_45 sn42_45 11.551961
Rsp41_46 sp41_46 sp42_46 11.551961
Rsn41_46 sn41_46 sn42_46 11.551961
Rsp41_47 sp41_47 sp42_47 11.551961
Rsn41_47 sn41_47 sn42_47 11.551961
Rsp41_48 sp41_48 sp42_48 11.551961
Rsn41_48 sn41_48 sn42_48 11.551961
Rsp41_49 sp41_49 sp42_49 11.551961
Rsn41_49 sn41_49 sn42_49 11.551961
Rsp41_50 sp41_50 sp42_50 11.551961
Rsn41_50 sn41_50 sn42_50 11.551961
Rsp41_51 sp41_51 sp42_51 11.551961
Rsn41_51 sn41_51 sn42_51 11.551961
Rsp41_52 sp41_52 sp42_52 11.551961
Rsn41_52 sn41_52 sn42_52 11.551961
Rsp41_53 sp41_53 sp42_53 11.551961
Rsn41_53 sn41_53 sn42_53 11.551961
Rsp41_54 sp41_54 sp42_54 11.551961
Rsn41_54 sn41_54 sn42_54 11.551961
Rsp41_55 sp41_55 sp42_55 11.551961
Rsn41_55 sn41_55 sn42_55 11.551961
Rsp41_56 sp41_56 sp42_56 11.551961
Rsn41_56 sn41_56 sn42_56 11.551961
Rsp41_57 sp41_57 sp42_57 11.551961
Rsn41_57 sn41_57 sn42_57 11.551961
Rsp41_58 sp41_58 sp42_58 11.551961
Rsn41_58 sn41_58 sn42_58 11.551961
Rsp41_59 sp41_59 sp42_59 11.551961
Rsn41_59 sn41_59 sn42_59 11.551961
Rsp41_60 sp41_60 sp42_60 11.551961
Rsn41_60 sn41_60 sn42_60 11.551961
Rsp41_61 sp41_61 sp42_61 11.551961
Rsn41_61 sn41_61 sn42_61 11.551961
Rsp41_62 sp41_62 sp42_62 11.551961
Rsn41_62 sn41_62 sn42_62 11.551961
Rsp41_63 sp41_63 sp42_63 11.551961
Rsn41_63 sn41_63 sn42_63 11.551961
Rsp41_64 sp41_64 sp42_64 11.551961
Rsn41_64 sn41_64 sn42_64 11.551961
Rsp41_65 sp41_65 sp42_65 11.551961
Rsn41_65 sn41_65 sn42_65 11.551961
Rsp41_66 sp41_66 sp42_66 11.551961
Rsn41_66 sn41_66 sn42_66 11.551961
Rsp41_67 sp41_67 sp42_67 11.551961
Rsn41_67 sn41_67 sn42_67 11.551961
Rsp41_68 sp41_68 sp42_68 11.551961
Rsn41_68 sn41_68 sn42_68 11.551961
Rsp41_69 sp41_69 sp42_69 11.551961
Rsn41_69 sn41_69 sn42_69 11.551961
Rsp41_70 sp41_70 sp42_70 11.551961
Rsn41_70 sn41_70 sn42_70 11.551961
Rsp41_71 sp41_71 sp42_71 11.551961
Rsn41_71 sn41_71 sn42_71 11.551961
Rsp41_72 sp41_72 sp42_72 11.551961
Rsn41_72 sn41_72 sn42_72 11.551961
Rsp41_73 sp41_73 sp42_73 11.551961
Rsn41_73 sn41_73 sn42_73 11.551961
Rsp41_74 sp41_74 sp42_74 11.551961
Rsn41_74 sn41_74 sn42_74 11.551961
Rsp41_75 sp41_75 sp42_75 11.551961
Rsn41_75 sn41_75 sn42_75 11.551961
Rsp41_76 sp41_76 sp42_76 11.551961
Rsn41_76 sn41_76 sn42_76 11.551961
Rsp41_77 sp41_77 sp42_77 11.551961
Rsn41_77 sn41_77 sn42_77 11.551961
Rsp41_78 sp41_78 sp42_78 11.551961
Rsn41_78 sn41_78 sn42_78 11.551961
Rsp41_79 sp41_79 sp42_79 11.551961
Rsn41_79 sn41_79 sn42_79 11.551961
Rsp41_80 sp41_80 sp42_80 11.551961
Rsn41_80 sn41_80 sn42_80 11.551961
Rsp41_81 sp41_81 sp42_81 11.551961
Rsn41_81 sn41_81 sn42_81 11.551961
Rsp41_82 sp41_82 sp42_82 11.551961
Rsn41_82 sn41_82 sn42_82 11.551961
Rsp41_83 sp41_83 sp42_83 11.551961
Rsn41_83 sn41_83 sn42_83 11.551961
Rsp41_84 sp41_84 sp42_84 11.551961
Rsn41_84 sn41_84 sn42_84 11.551961
Rsp42_1 sp42_1 sp43_1 11.551961
Rsn42_1 sn42_1 sn43_1 11.551961
Rsp42_2 sp42_2 sp43_2 11.551961
Rsn42_2 sn42_2 sn43_2 11.551961
Rsp42_3 sp42_3 sp43_3 11.551961
Rsn42_3 sn42_3 sn43_3 11.551961
Rsp42_4 sp42_4 sp43_4 11.551961
Rsn42_4 sn42_4 sn43_4 11.551961
Rsp42_5 sp42_5 sp43_5 11.551961
Rsn42_5 sn42_5 sn43_5 11.551961
Rsp42_6 sp42_6 sp43_6 11.551961
Rsn42_6 sn42_6 sn43_6 11.551961
Rsp42_7 sp42_7 sp43_7 11.551961
Rsn42_7 sn42_7 sn43_7 11.551961
Rsp42_8 sp42_8 sp43_8 11.551961
Rsn42_8 sn42_8 sn43_8 11.551961
Rsp42_9 sp42_9 sp43_9 11.551961
Rsn42_9 sn42_9 sn43_9 11.551961
Rsp42_10 sp42_10 sp43_10 11.551961
Rsn42_10 sn42_10 sn43_10 11.551961
Rsp42_11 sp42_11 sp43_11 11.551961
Rsn42_11 sn42_11 sn43_11 11.551961
Rsp42_12 sp42_12 sp43_12 11.551961
Rsn42_12 sn42_12 sn43_12 11.551961
Rsp42_13 sp42_13 sp43_13 11.551961
Rsn42_13 sn42_13 sn43_13 11.551961
Rsp42_14 sp42_14 sp43_14 11.551961
Rsn42_14 sn42_14 sn43_14 11.551961
Rsp42_15 sp42_15 sp43_15 11.551961
Rsn42_15 sn42_15 sn43_15 11.551961
Rsp42_16 sp42_16 sp43_16 11.551961
Rsn42_16 sn42_16 sn43_16 11.551961
Rsp42_17 sp42_17 sp43_17 11.551961
Rsn42_17 sn42_17 sn43_17 11.551961
Rsp42_18 sp42_18 sp43_18 11.551961
Rsn42_18 sn42_18 sn43_18 11.551961
Rsp42_19 sp42_19 sp43_19 11.551961
Rsn42_19 sn42_19 sn43_19 11.551961
Rsp42_20 sp42_20 sp43_20 11.551961
Rsn42_20 sn42_20 sn43_20 11.551961
Rsp42_21 sp42_21 sp43_21 11.551961
Rsn42_21 sn42_21 sn43_21 11.551961
Rsp42_22 sp42_22 sp43_22 11.551961
Rsn42_22 sn42_22 sn43_22 11.551961
Rsp42_23 sp42_23 sp43_23 11.551961
Rsn42_23 sn42_23 sn43_23 11.551961
Rsp42_24 sp42_24 sp43_24 11.551961
Rsn42_24 sn42_24 sn43_24 11.551961
Rsp42_25 sp42_25 sp43_25 11.551961
Rsn42_25 sn42_25 sn43_25 11.551961
Rsp42_26 sp42_26 sp43_26 11.551961
Rsn42_26 sn42_26 sn43_26 11.551961
Rsp42_27 sp42_27 sp43_27 11.551961
Rsn42_27 sn42_27 sn43_27 11.551961
Rsp42_28 sp42_28 sp43_28 11.551961
Rsn42_28 sn42_28 sn43_28 11.551961
Rsp42_29 sp42_29 sp43_29 11.551961
Rsn42_29 sn42_29 sn43_29 11.551961
Rsp42_30 sp42_30 sp43_30 11.551961
Rsn42_30 sn42_30 sn43_30 11.551961
Rsp42_31 sp42_31 sp43_31 11.551961
Rsn42_31 sn42_31 sn43_31 11.551961
Rsp42_32 sp42_32 sp43_32 11.551961
Rsn42_32 sn42_32 sn43_32 11.551961
Rsp42_33 sp42_33 sp43_33 11.551961
Rsn42_33 sn42_33 sn43_33 11.551961
Rsp42_34 sp42_34 sp43_34 11.551961
Rsn42_34 sn42_34 sn43_34 11.551961
Rsp42_35 sp42_35 sp43_35 11.551961
Rsn42_35 sn42_35 sn43_35 11.551961
Rsp42_36 sp42_36 sp43_36 11.551961
Rsn42_36 sn42_36 sn43_36 11.551961
Rsp42_37 sp42_37 sp43_37 11.551961
Rsn42_37 sn42_37 sn43_37 11.551961
Rsp42_38 sp42_38 sp43_38 11.551961
Rsn42_38 sn42_38 sn43_38 11.551961
Rsp42_39 sp42_39 sp43_39 11.551961
Rsn42_39 sn42_39 sn43_39 11.551961
Rsp42_40 sp42_40 sp43_40 11.551961
Rsn42_40 sn42_40 sn43_40 11.551961
Rsp42_41 sp42_41 sp43_41 11.551961
Rsn42_41 sn42_41 sn43_41 11.551961
Rsp42_42 sp42_42 sp43_42 11.551961
Rsn42_42 sn42_42 sn43_42 11.551961
Rsp42_43 sp42_43 sp43_43 11.551961
Rsn42_43 sn42_43 sn43_43 11.551961
Rsp42_44 sp42_44 sp43_44 11.551961
Rsn42_44 sn42_44 sn43_44 11.551961
Rsp42_45 sp42_45 sp43_45 11.551961
Rsn42_45 sn42_45 sn43_45 11.551961
Rsp42_46 sp42_46 sp43_46 11.551961
Rsn42_46 sn42_46 sn43_46 11.551961
Rsp42_47 sp42_47 sp43_47 11.551961
Rsn42_47 sn42_47 sn43_47 11.551961
Rsp42_48 sp42_48 sp43_48 11.551961
Rsn42_48 sn42_48 sn43_48 11.551961
Rsp42_49 sp42_49 sp43_49 11.551961
Rsn42_49 sn42_49 sn43_49 11.551961
Rsp42_50 sp42_50 sp43_50 11.551961
Rsn42_50 sn42_50 sn43_50 11.551961
Rsp42_51 sp42_51 sp43_51 11.551961
Rsn42_51 sn42_51 sn43_51 11.551961
Rsp42_52 sp42_52 sp43_52 11.551961
Rsn42_52 sn42_52 sn43_52 11.551961
Rsp42_53 sp42_53 sp43_53 11.551961
Rsn42_53 sn42_53 sn43_53 11.551961
Rsp42_54 sp42_54 sp43_54 11.551961
Rsn42_54 sn42_54 sn43_54 11.551961
Rsp42_55 sp42_55 sp43_55 11.551961
Rsn42_55 sn42_55 sn43_55 11.551961
Rsp42_56 sp42_56 sp43_56 11.551961
Rsn42_56 sn42_56 sn43_56 11.551961
Rsp42_57 sp42_57 sp43_57 11.551961
Rsn42_57 sn42_57 sn43_57 11.551961
Rsp42_58 sp42_58 sp43_58 11.551961
Rsn42_58 sn42_58 sn43_58 11.551961
Rsp42_59 sp42_59 sp43_59 11.551961
Rsn42_59 sn42_59 sn43_59 11.551961
Rsp42_60 sp42_60 sp43_60 11.551961
Rsn42_60 sn42_60 sn43_60 11.551961
Rsp42_61 sp42_61 sp43_61 11.551961
Rsn42_61 sn42_61 sn43_61 11.551961
Rsp42_62 sp42_62 sp43_62 11.551961
Rsn42_62 sn42_62 sn43_62 11.551961
Rsp42_63 sp42_63 sp43_63 11.551961
Rsn42_63 sn42_63 sn43_63 11.551961
Rsp42_64 sp42_64 sp43_64 11.551961
Rsn42_64 sn42_64 sn43_64 11.551961
Rsp42_65 sp42_65 sp43_65 11.551961
Rsn42_65 sn42_65 sn43_65 11.551961
Rsp42_66 sp42_66 sp43_66 11.551961
Rsn42_66 sn42_66 sn43_66 11.551961
Rsp42_67 sp42_67 sp43_67 11.551961
Rsn42_67 sn42_67 sn43_67 11.551961
Rsp42_68 sp42_68 sp43_68 11.551961
Rsn42_68 sn42_68 sn43_68 11.551961
Rsp42_69 sp42_69 sp43_69 11.551961
Rsn42_69 sn42_69 sn43_69 11.551961
Rsp42_70 sp42_70 sp43_70 11.551961
Rsn42_70 sn42_70 sn43_70 11.551961
Rsp42_71 sp42_71 sp43_71 11.551961
Rsn42_71 sn42_71 sn43_71 11.551961
Rsp42_72 sp42_72 sp43_72 11.551961
Rsn42_72 sn42_72 sn43_72 11.551961
Rsp42_73 sp42_73 sp43_73 11.551961
Rsn42_73 sn42_73 sn43_73 11.551961
Rsp42_74 sp42_74 sp43_74 11.551961
Rsn42_74 sn42_74 sn43_74 11.551961
Rsp42_75 sp42_75 sp43_75 11.551961
Rsn42_75 sn42_75 sn43_75 11.551961
Rsp42_76 sp42_76 sp43_76 11.551961
Rsn42_76 sn42_76 sn43_76 11.551961
Rsp42_77 sp42_77 sp43_77 11.551961
Rsn42_77 sn42_77 sn43_77 11.551961
Rsp42_78 sp42_78 sp43_78 11.551961
Rsn42_78 sn42_78 sn43_78 11.551961
Rsp42_79 sp42_79 sp43_79 11.551961
Rsn42_79 sn42_79 sn43_79 11.551961
Rsp42_80 sp42_80 sp43_80 11.551961
Rsn42_80 sn42_80 sn43_80 11.551961
Rsp42_81 sp42_81 sp43_81 11.551961
Rsn42_81 sn42_81 sn43_81 11.551961
Rsp42_82 sp42_82 sp43_82 11.551961
Rsn42_82 sn42_82 sn43_82 11.551961
Rsp42_83 sp42_83 sp43_83 11.551961
Rsn42_83 sn42_83 sn43_83 11.551961
Rsp42_84 sp42_84 sp43_84 11.551961
Rsn42_84 sn42_84 sn43_84 11.551961
Rsp43_1 sp43_1 sp44_1 11.551961
Rsn43_1 sn43_1 sn44_1 11.551961
Rsp43_2 sp43_2 sp44_2 11.551961
Rsn43_2 sn43_2 sn44_2 11.551961
Rsp43_3 sp43_3 sp44_3 11.551961
Rsn43_3 sn43_3 sn44_3 11.551961
Rsp43_4 sp43_4 sp44_4 11.551961
Rsn43_4 sn43_4 sn44_4 11.551961
Rsp43_5 sp43_5 sp44_5 11.551961
Rsn43_5 sn43_5 sn44_5 11.551961
Rsp43_6 sp43_6 sp44_6 11.551961
Rsn43_6 sn43_6 sn44_6 11.551961
Rsp43_7 sp43_7 sp44_7 11.551961
Rsn43_7 sn43_7 sn44_7 11.551961
Rsp43_8 sp43_8 sp44_8 11.551961
Rsn43_8 sn43_8 sn44_8 11.551961
Rsp43_9 sp43_9 sp44_9 11.551961
Rsn43_9 sn43_9 sn44_9 11.551961
Rsp43_10 sp43_10 sp44_10 11.551961
Rsn43_10 sn43_10 sn44_10 11.551961
Rsp43_11 sp43_11 sp44_11 11.551961
Rsn43_11 sn43_11 sn44_11 11.551961
Rsp43_12 sp43_12 sp44_12 11.551961
Rsn43_12 sn43_12 sn44_12 11.551961
Rsp43_13 sp43_13 sp44_13 11.551961
Rsn43_13 sn43_13 sn44_13 11.551961
Rsp43_14 sp43_14 sp44_14 11.551961
Rsn43_14 sn43_14 sn44_14 11.551961
Rsp43_15 sp43_15 sp44_15 11.551961
Rsn43_15 sn43_15 sn44_15 11.551961
Rsp43_16 sp43_16 sp44_16 11.551961
Rsn43_16 sn43_16 sn44_16 11.551961
Rsp43_17 sp43_17 sp44_17 11.551961
Rsn43_17 sn43_17 sn44_17 11.551961
Rsp43_18 sp43_18 sp44_18 11.551961
Rsn43_18 sn43_18 sn44_18 11.551961
Rsp43_19 sp43_19 sp44_19 11.551961
Rsn43_19 sn43_19 sn44_19 11.551961
Rsp43_20 sp43_20 sp44_20 11.551961
Rsn43_20 sn43_20 sn44_20 11.551961
Rsp43_21 sp43_21 sp44_21 11.551961
Rsn43_21 sn43_21 sn44_21 11.551961
Rsp43_22 sp43_22 sp44_22 11.551961
Rsn43_22 sn43_22 sn44_22 11.551961
Rsp43_23 sp43_23 sp44_23 11.551961
Rsn43_23 sn43_23 sn44_23 11.551961
Rsp43_24 sp43_24 sp44_24 11.551961
Rsn43_24 sn43_24 sn44_24 11.551961
Rsp43_25 sp43_25 sp44_25 11.551961
Rsn43_25 sn43_25 sn44_25 11.551961
Rsp43_26 sp43_26 sp44_26 11.551961
Rsn43_26 sn43_26 sn44_26 11.551961
Rsp43_27 sp43_27 sp44_27 11.551961
Rsn43_27 sn43_27 sn44_27 11.551961
Rsp43_28 sp43_28 sp44_28 11.551961
Rsn43_28 sn43_28 sn44_28 11.551961
Rsp43_29 sp43_29 sp44_29 11.551961
Rsn43_29 sn43_29 sn44_29 11.551961
Rsp43_30 sp43_30 sp44_30 11.551961
Rsn43_30 sn43_30 sn44_30 11.551961
Rsp43_31 sp43_31 sp44_31 11.551961
Rsn43_31 sn43_31 sn44_31 11.551961
Rsp43_32 sp43_32 sp44_32 11.551961
Rsn43_32 sn43_32 sn44_32 11.551961
Rsp43_33 sp43_33 sp44_33 11.551961
Rsn43_33 sn43_33 sn44_33 11.551961
Rsp43_34 sp43_34 sp44_34 11.551961
Rsn43_34 sn43_34 sn44_34 11.551961
Rsp43_35 sp43_35 sp44_35 11.551961
Rsn43_35 sn43_35 sn44_35 11.551961
Rsp43_36 sp43_36 sp44_36 11.551961
Rsn43_36 sn43_36 sn44_36 11.551961
Rsp43_37 sp43_37 sp44_37 11.551961
Rsn43_37 sn43_37 sn44_37 11.551961
Rsp43_38 sp43_38 sp44_38 11.551961
Rsn43_38 sn43_38 sn44_38 11.551961
Rsp43_39 sp43_39 sp44_39 11.551961
Rsn43_39 sn43_39 sn44_39 11.551961
Rsp43_40 sp43_40 sp44_40 11.551961
Rsn43_40 sn43_40 sn44_40 11.551961
Rsp43_41 sp43_41 sp44_41 11.551961
Rsn43_41 sn43_41 sn44_41 11.551961
Rsp43_42 sp43_42 sp44_42 11.551961
Rsn43_42 sn43_42 sn44_42 11.551961
Rsp43_43 sp43_43 sp44_43 11.551961
Rsn43_43 sn43_43 sn44_43 11.551961
Rsp43_44 sp43_44 sp44_44 11.551961
Rsn43_44 sn43_44 sn44_44 11.551961
Rsp43_45 sp43_45 sp44_45 11.551961
Rsn43_45 sn43_45 sn44_45 11.551961
Rsp43_46 sp43_46 sp44_46 11.551961
Rsn43_46 sn43_46 sn44_46 11.551961
Rsp43_47 sp43_47 sp44_47 11.551961
Rsn43_47 sn43_47 sn44_47 11.551961
Rsp43_48 sp43_48 sp44_48 11.551961
Rsn43_48 sn43_48 sn44_48 11.551961
Rsp43_49 sp43_49 sp44_49 11.551961
Rsn43_49 sn43_49 sn44_49 11.551961
Rsp43_50 sp43_50 sp44_50 11.551961
Rsn43_50 sn43_50 sn44_50 11.551961
Rsp43_51 sp43_51 sp44_51 11.551961
Rsn43_51 sn43_51 sn44_51 11.551961
Rsp43_52 sp43_52 sp44_52 11.551961
Rsn43_52 sn43_52 sn44_52 11.551961
Rsp43_53 sp43_53 sp44_53 11.551961
Rsn43_53 sn43_53 sn44_53 11.551961
Rsp43_54 sp43_54 sp44_54 11.551961
Rsn43_54 sn43_54 sn44_54 11.551961
Rsp43_55 sp43_55 sp44_55 11.551961
Rsn43_55 sn43_55 sn44_55 11.551961
Rsp43_56 sp43_56 sp44_56 11.551961
Rsn43_56 sn43_56 sn44_56 11.551961
Rsp43_57 sp43_57 sp44_57 11.551961
Rsn43_57 sn43_57 sn44_57 11.551961
Rsp43_58 sp43_58 sp44_58 11.551961
Rsn43_58 sn43_58 sn44_58 11.551961
Rsp43_59 sp43_59 sp44_59 11.551961
Rsn43_59 sn43_59 sn44_59 11.551961
Rsp43_60 sp43_60 sp44_60 11.551961
Rsn43_60 sn43_60 sn44_60 11.551961
Rsp43_61 sp43_61 sp44_61 11.551961
Rsn43_61 sn43_61 sn44_61 11.551961
Rsp43_62 sp43_62 sp44_62 11.551961
Rsn43_62 sn43_62 sn44_62 11.551961
Rsp43_63 sp43_63 sp44_63 11.551961
Rsn43_63 sn43_63 sn44_63 11.551961
Rsp43_64 sp43_64 sp44_64 11.551961
Rsn43_64 sn43_64 sn44_64 11.551961
Rsp43_65 sp43_65 sp44_65 11.551961
Rsn43_65 sn43_65 sn44_65 11.551961
Rsp43_66 sp43_66 sp44_66 11.551961
Rsn43_66 sn43_66 sn44_66 11.551961
Rsp43_67 sp43_67 sp44_67 11.551961
Rsn43_67 sn43_67 sn44_67 11.551961
Rsp43_68 sp43_68 sp44_68 11.551961
Rsn43_68 sn43_68 sn44_68 11.551961
Rsp43_69 sp43_69 sp44_69 11.551961
Rsn43_69 sn43_69 sn44_69 11.551961
Rsp43_70 sp43_70 sp44_70 11.551961
Rsn43_70 sn43_70 sn44_70 11.551961
Rsp43_71 sp43_71 sp44_71 11.551961
Rsn43_71 sn43_71 sn44_71 11.551961
Rsp43_72 sp43_72 sp44_72 11.551961
Rsn43_72 sn43_72 sn44_72 11.551961
Rsp43_73 sp43_73 sp44_73 11.551961
Rsn43_73 sn43_73 sn44_73 11.551961
Rsp43_74 sp43_74 sp44_74 11.551961
Rsn43_74 sn43_74 sn44_74 11.551961
Rsp43_75 sp43_75 sp44_75 11.551961
Rsn43_75 sn43_75 sn44_75 11.551961
Rsp43_76 sp43_76 sp44_76 11.551961
Rsn43_76 sn43_76 sn44_76 11.551961
Rsp43_77 sp43_77 sp44_77 11.551961
Rsn43_77 sn43_77 sn44_77 11.551961
Rsp43_78 sp43_78 sp44_78 11.551961
Rsn43_78 sn43_78 sn44_78 11.551961
Rsp43_79 sp43_79 sp44_79 11.551961
Rsn43_79 sn43_79 sn44_79 11.551961
Rsp43_80 sp43_80 sp44_80 11.551961
Rsn43_80 sn43_80 sn44_80 11.551961
Rsp43_81 sp43_81 sp44_81 11.551961
Rsn43_81 sn43_81 sn44_81 11.551961
Rsp43_82 sp43_82 sp44_82 11.551961
Rsn43_82 sn43_82 sn44_82 11.551961
Rsp43_83 sp43_83 sp44_83 11.551961
Rsn43_83 sn43_83 sn44_83 11.551961
Rsp43_84 sp43_84 sp44_84 11.551961
Rsn43_84 sn43_84 sn44_84 11.551961
Rsp44_1 sp44_1 sp45_1 11.551961
Rsn44_1 sn44_1 sn45_1 11.551961
Rsp44_2 sp44_2 sp45_2 11.551961
Rsn44_2 sn44_2 sn45_2 11.551961
Rsp44_3 sp44_3 sp45_3 11.551961
Rsn44_3 sn44_3 sn45_3 11.551961
Rsp44_4 sp44_4 sp45_4 11.551961
Rsn44_4 sn44_4 sn45_4 11.551961
Rsp44_5 sp44_5 sp45_5 11.551961
Rsn44_5 sn44_5 sn45_5 11.551961
Rsp44_6 sp44_6 sp45_6 11.551961
Rsn44_6 sn44_6 sn45_6 11.551961
Rsp44_7 sp44_7 sp45_7 11.551961
Rsn44_7 sn44_7 sn45_7 11.551961
Rsp44_8 sp44_8 sp45_8 11.551961
Rsn44_8 sn44_8 sn45_8 11.551961
Rsp44_9 sp44_9 sp45_9 11.551961
Rsn44_9 sn44_9 sn45_9 11.551961
Rsp44_10 sp44_10 sp45_10 11.551961
Rsn44_10 sn44_10 sn45_10 11.551961
Rsp44_11 sp44_11 sp45_11 11.551961
Rsn44_11 sn44_11 sn45_11 11.551961
Rsp44_12 sp44_12 sp45_12 11.551961
Rsn44_12 sn44_12 sn45_12 11.551961
Rsp44_13 sp44_13 sp45_13 11.551961
Rsn44_13 sn44_13 sn45_13 11.551961
Rsp44_14 sp44_14 sp45_14 11.551961
Rsn44_14 sn44_14 sn45_14 11.551961
Rsp44_15 sp44_15 sp45_15 11.551961
Rsn44_15 sn44_15 sn45_15 11.551961
Rsp44_16 sp44_16 sp45_16 11.551961
Rsn44_16 sn44_16 sn45_16 11.551961
Rsp44_17 sp44_17 sp45_17 11.551961
Rsn44_17 sn44_17 sn45_17 11.551961
Rsp44_18 sp44_18 sp45_18 11.551961
Rsn44_18 sn44_18 sn45_18 11.551961
Rsp44_19 sp44_19 sp45_19 11.551961
Rsn44_19 sn44_19 sn45_19 11.551961
Rsp44_20 sp44_20 sp45_20 11.551961
Rsn44_20 sn44_20 sn45_20 11.551961
Rsp44_21 sp44_21 sp45_21 11.551961
Rsn44_21 sn44_21 sn45_21 11.551961
Rsp44_22 sp44_22 sp45_22 11.551961
Rsn44_22 sn44_22 sn45_22 11.551961
Rsp44_23 sp44_23 sp45_23 11.551961
Rsn44_23 sn44_23 sn45_23 11.551961
Rsp44_24 sp44_24 sp45_24 11.551961
Rsn44_24 sn44_24 sn45_24 11.551961
Rsp44_25 sp44_25 sp45_25 11.551961
Rsn44_25 sn44_25 sn45_25 11.551961
Rsp44_26 sp44_26 sp45_26 11.551961
Rsn44_26 sn44_26 sn45_26 11.551961
Rsp44_27 sp44_27 sp45_27 11.551961
Rsn44_27 sn44_27 sn45_27 11.551961
Rsp44_28 sp44_28 sp45_28 11.551961
Rsn44_28 sn44_28 sn45_28 11.551961
Rsp44_29 sp44_29 sp45_29 11.551961
Rsn44_29 sn44_29 sn45_29 11.551961
Rsp44_30 sp44_30 sp45_30 11.551961
Rsn44_30 sn44_30 sn45_30 11.551961
Rsp44_31 sp44_31 sp45_31 11.551961
Rsn44_31 sn44_31 sn45_31 11.551961
Rsp44_32 sp44_32 sp45_32 11.551961
Rsn44_32 sn44_32 sn45_32 11.551961
Rsp44_33 sp44_33 sp45_33 11.551961
Rsn44_33 sn44_33 sn45_33 11.551961
Rsp44_34 sp44_34 sp45_34 11.551961
Rsn44_34 sn44_34 sn45_34 11.551961
Rsp44_35 sp44_35 sp45_35 11.551961
Rsn44_35 sn44_35 sn45_35 11.551961
Rsp44_36 sp44_36 sp45_36 11.551961
Rsn44_36 sn44_36 sn45_36 11.551961
Rsp44_37 sp44_37 sp45_37 11.551961
Rsn44_37 sn44_37 sn45_37 11.551961
Rsp44_38 sp44_38 sp45_38 11.551961
Rsn44_38 sn44_38 sn45_38 11.551961
Rsp44_39 sp44_39 sp45_39 11.551961
Rsn44_39 sn44_39 sn45_39 11.551961
Rsp44_40 sp44_40 sp45_40 11.551961
Rsn44_40 sn44_40 sn45_40 11.551961
Rsp44_41 sp44_41 sp45_41 11.551961
Rsn44_41 sn44_41 sn45_41 11.551961
Rsp44_42 sp44_42 sp45_42 11.551961
Rsn44_42 sn44_42 sn45_42 11.551961
Rsp44_43 sp44_43 sp45_43 11.551961
Rsn44_43 sn44_43 sn45_43 11.551961
Rsp44_44 sp44_44 sp45_44 11.551961
Rsn44_44 sn44_44 sn45_44 11.551961
Rsp44_45 sp44_45 sp45_45 11.551961
Rsn44_45 sn44_45 sn45_45 11.551961
Rsp44_46 sp44_46 sp45_46 11.551961
Rsn44_46 sn44_46 sn45_46 11.551961
Rsp44_47 sp44_47 sp45_47 11.551961
Rsn44_47 sn44_47 sn45_47 11.551961
Rsp44_48 sp44_48 sp45_48 11.551961
Rsn44_48 sn44_48 sn45_48 11.551961
Rsp44_49 sp44_49 sp45_49 11.551961
Rsn44_49 sn44_49 sn45_49 11.551961
Rsp44_50 sp44_50 sp45_50 11.551961
Rsn44_50 sn44_50 sn45_50 11.551961
Rsp44_51 sp44_51 sp45_51 11.551961
Rsn44_51 sn44_51 sn45_51 11.551961
Rsp44_52 sp44_52 sp45_52 11.551961
Rsn44_52 sn44_52 sn45_52 11.551961
Rsp44_53 sp44_53 sp45_53 11.551961
Rsn44_53 sn44_53 sn45_53 11.551961
Rsp44_54 sp44_54 sp45_54 11.551961
Rsn44_54 sn44_54 sn45_54 11.551961
Rsp44_55 sp44_55 sp45_55 11.551961
Rsn44_55 sn44_55 sn45_55 11.551961
Rsp44_56 sp44_56 sp45_56 11.551961
Rsn44_56 sn44_56 sn45_56 11.551961
Rsp44_57 sp44_57 sp45_57 11.551961
Rsn44_57 sn44_57 sn45_57 11.551961
Rsp44_58 sp44_58 sp45_58 11.551961
Rsn44_58 sn44_58 sn45_58 11.551961
Rsp44_59 sp44_59 sp45_59 11.551961
Rsn44_59 sn44_59 sn45_59 11.551961
Rsp44_60 sp44_60 sp45_60 11.551961
Rsn44_60 sn44_60 sn45_60 11.551961
Rsp44_61 sp44_61 sp45_61 11.551961
Rsn44_61 sn44_61 sn45_61 11.551961
Rsp44_62 sp44_62 sp45_62 11.551961
Rsn44_62 sn44_62 sn45_62 11.551961
Rsp44_63 sp44_63 sp45_63 11.551961
Rsn44_63 sn44_63 sn45_63 11.551961
Rsp44_64 sp44_64 sp45_64 11.551961
Rsn44_64 sn44_64 sn45_64 11.551961
Rsp44_65 sp44_65 sp45_65 11.551961
Rsn44_65 sn44_65 sn45_65 11.551961
Rsp44_66 sp44_66 sp45_66 11.551961
Rsn44_66 sn44_66 sn45_66 11.551961
Rsp44_67 sp44_67 sp45_67 11.551961
Rsn44_67 sn44_67 sn45_67 11.551961
Rsp44_68 sp44_68 sp45_68 11.551961
Rsn44_68 sn44_68 sn45_68 11.551961
Rsp44_69 sp44_69 sp45_69 11.551961
Rsn44_69 sn44_69 sn45_69 11.551961
Rsp44_70 sp44_70 sp45_70 11.551961
Rsn44_70 sn44_70 sn45_70 11.551961
Rsp44_71 sp44_71 sp45_71 11.551961
Rsn44_71 sn44_71 sn45_71 11.551961
Rsp44_72 sp44_72 sp45_72 11.551961
Rsn44_72 sn44_72 sn45_72 11.551961
Rsp44_73 sp44_73 sp45_73 11.551961
Rsn44_73 sn44_73 sn45_73 11.551961
Rsp44_74 sp44_74 sp45_74 11.551961
Rsn44_74 sn44_74 sn45_74 11.551961
Rsp44_75 sp44_75 sp45_75 11.551961
Rsn44_75 sn44_75 sn45_75 11.551961
Rsp44_76 sp44_76 sp45_76 11.551961
Rsn44_76 sn44_76 sn45_76 11.551961
Rsp44_77 sp44_77 sp45_77 11.551961
Rsn44_77 sn44_77 sn45_77 11.551961
Rsp44_78 sp44_78 sp45_78 11.551961
Rsn44_78 sn44_78 sn45_78 11.551961
Rsp44_79 sp44_79 sp45_79 11.551961
Rsn44_79 sn44_79 sn45_79 11.551961
Rsp44_80 sp44_80 sp45_80 11.551961
Rsn44_80 sn44_80 sn45_80 11.551961
Rsp44_81 sp44_81 sp45_81 11.551961
Rsn44_81 sn44_81 sn45_81 11.551961
Rsp44_82 sp44_82 sp45_82 11.551961
Rsn44_82 sn44_82 sn45_82 11.551961
Rsp44_83 sp44_83 sp45_83 11.551961
Rsn44_83 sn44_83 sn45_83 11.551961
Rsp44_84 sp44_84 sp45_84 11.551961
Rsn44_84 sn44_84 sn45_84 11.551961
Rsp45_1 sp45_1 sp46_1 11.551961
Rsn45_1 sn45_1 sn46_1 11.551961
Rsp45_2 sp45_2 sp46_2 11.551961
Rsn45_2 sn45_2 sn46_2 11.551961
Rsp45_3 sp45_3 sp46_3 11.551961
Rsn45_3 sn45_3 sn46_3 11.551961
Rsp45_4 sp45_4 sp46_4 11.551961
Rsn45_4 sn45_4 sn46_4 11.551961
Rsp45_5 sp45_5 sp46_5 11.551961
Rsn45_5 sn45_5 sn46_5 11.551961
Rsp45_6 sp45_6 sp46_6 11.551961
Rsn45_6 sn45_6 sn46_6 11.551961
Rsp45_7 sp45_7 sp46_7 11.551961
Rsn45_7 sn45_7 sn46_7 11.551961
Rsp45_8 sp45_8 sp46_8 11.551961
Rsn45_8 sn45_8 sn46_8 11.551961
Rsp45_9 sp45_9 sp46_9 11.551961
Rsn45_9 sn45_9 sn46_9 11.551961
Rsp45_10 sp45_10 sp46_10 11.551961
Rsn45_10 sn45_10 sn46_10 11.551961
Rsp45_11 sp45_11 sp46_11 11.551961
Rsn45_11 sn45_11 sn46_11 11.551961
Rsp45_12 sp45_12 sp46_12 11.551961
Rsn45_12 sn45_12 sn46_12 11.551961
Rsp45_13 sp45_13 sp46_13 11.551961
Rsn45_13 sn45_13 sn46_13 11.551961
Rsp45_14 sp45_14 sp46_14 11.551961
Rsn45_14 sn45_14 sn46_14 11.551961
Rsp45_15 sp45_15 sp46_15 11.551961
Rsn45_15 sn45_15 sn46_15 11.551961
Rsp45_16 sp45_16 sp46_16 11.551961
Rsn45_16 sn45_16 sn46_16 11.551961
Rsp45_17 sp45_17 sp46_17 11.551961
Rsn45_17 sn45_17 sn46_17 11.551961
Rsp45_18 sp45_18 sp46_18 11.551961
Rsn45_18 sn45_18 sn46_18 11.551961
Rsp45_19 sp45_19 sp46_19 11.551961
Rsn45_19 sn45_19 sn46_19 11.551961
Rsp45_20 sp45_20 sp46_20 11.551961
Rsn45_20 sn45_20 sn46_20 11.551961
Rsp45_21 sp45_21 sp46_21 11.551961
Rsn45_21 sn45_21 sn46_21 11.551961
Rsp45_22 sp45_22 sp46_22 11.551961
Rsn45_22 sn45_22 sn46_22 11.551961
Rsp45_23 sp45_23 sp46_23 11.551961
Rsn45_23 sn45_23 sn46_23 11.551961
Rsp45_24 sp45_24 sp46_24 11.551961
Rsn45_24 sn45_24 sn46_24 11.551961
Rsp45_25 sp45_25 sp46_25 11.551961
Rsn45_25 sn45_25 sn46_25 11.551961
Rsp45_26 sp45_26 sp46_26 11.551961
Rsn45_26 sn45_26 sn46_26 11.551961
Rsp45_27 sp45_27 sp46_27 11.551961
Rsn45_27 sn45_27 sn46_27 11.551961
Rsp45_28 sp45_28 sp46_28 11.551961
Rsn45_28 sn45_28 sn46_28 11.551961
Rsp45_29 sp45_29 sp46_29 11.551961
Rsn45_29 sn45_29 sn46_29 11.551961
Rsp45_30 sp45_30 sp46_30 11.551961
Rsn45_30 sn45_30 sn46_30 11.551961
Rsp45_31 sp45_31 sp46_31 11.551961
Rsn45_31 sn45_31 sn46_31 11.551961
Rsp45_32 sp45_32 sp46_32 11.551961
Rsn45_32 sn45_32 sn46_32 11.551961
Rsp45_33 sp45_33 sp46_33 11.551961
Rsn45_33 sn45_33 sn46_33 11.551961
Rsp45_34 sp45_34 sp46_34 11.551961
Rsn45_34 sn45_34 sn46_34 11.551961
Rsp45_35 sp45_35 sp46_35 11.551961
Rsn45_35 sn45_35 sn46_35 11.551961
Rsp45_36 sp45_36 sp46_36 11.551961
Rsn45_36 sn45_36 sn46_36 11.551961
Rsp45_37 sp45_37 sp46_37 11.551961
Rsn45_37 sn45_37 sn46_37 11.551961
Rsp45_38 sp45_38 sp46_38 11.551961
Rsn45_38 sn45_38 sn46_38 11.551961
Rsp45_39 sp45_39 sp46_39 11.551961
Rsn45_39 sn45_39 sn46_39 11.551961
Rsp45_40 sp45_40 sp46_40 11.551961
Rsn45_40 sn45_40 sn46_40 11.551961
Rsp45_41 sp45_41 sp46_41 11.551961
Rsn45_41 sn45_41 sn46_41 11.551961
Rsp45_42 sp45_42 sp46_42 11.551961
Rsn45_42 sn45_42 sn46_42 11.551961
Rsp45_43 sp45_43 sp46_43 11.551961
Rsn45_43 sn45_43 sn46_43 11.551961
Rsp45_44 sp45_44 sp46_44 11.551961
Rsn45_44 sn45_44 sn46_44 11.551961
Rsp45_45 sp45_45 sp46_45 11.551961
Rsn45_45 sn45_45 sn46_45 11.551961
Rsp45_46 sp45_46 sp46_46 11.551961
Rsn45_46 sn45_46 sn46_46 11.551961
Rsp45_47 sp45_47 sp46_47 11.551961
Rsn45_47 sn45_47 sn46_47 11.551961
Rsp45_48 sp45_48 sp46_48 11.551961
Rsn45_48 sn45_48 sn46_48 11.551961
Rsp45_49 sp45_49 sp46_49 11.551961
Rsn45_49 sn45_49 sn46_49 11.551961
Rsp45_50 sp45_50 sp46_50 11.551961
Rsn45_50 sn45_50 sn46_50 11.551961
Rsp45_51 sp45_51 sp46_51 11.551961
Rsn45_51 sn45_51 sn46_51 11.551961
Rsp45_52 sp45_52 sp46_52 11.551961
Rsn45_52 sn45_52 sn46_52 11.551961
Rsp45_53 sp45_53 sp46_53 11.551961
Rsn45_53 sn45_53 sn46_53 11.551961
Rsp45_54 sp45_54 sp46_54 11.551961
Rsn45_54 sn45_54 sn46_54 11.551961
Rsp45_55 sp45_55 sp46_55 11.551961
Rsn45_55 sn45_55 sn46_55 11.551961
Rsp45_56 sp45_56 sp46_56 11.551961
Rsn45_56 sn45_56 sn46_56 11.551961
Rsp45_57 sp45_57 sp46_57 11.551961
Rsn45_57 sn45_57 sn46_57 11.551961
Rsp45_58 sp45_58 sp46_58 11.551961
Rsn45_58 sn45_58 sn46_58 11.551961
Rsp45_59 sp45_59 sp46_59 11.551961
Rsn45_59 sn45_59 sn46_59 11.551961
Rsp45_60 sp45_60 sp46_60 11.551961
Rsn45_60 sn45_60 sn46_60 11.551961
Rsp45_61 sp45_61 sp46_61 11.551961
Rsn45_61 sn45_61 sn46_61 11.551961
Rsp45_62 sp45_62 sp46_62 11.551961
Rsn45_62 sn45_62 sn46_62 11.551961
Rsp45_63 sp45_63 sp46_63 11.551961
Rsn45_63 sn45_63 sn46_63 11.551961
Rsp45_64 sp45_64 sp46_64 11.551961
Rsn45_64 sn45_64 sn46_64 11.551961
Rsp45_65 sp45_65 sp46_65 11.551961
Rsn45_65 sn45_65 sn46_65 11.551961
Rsp45_66 sp45_66 sp46_66 11.551961
Rsn45_66 sn45_66 sn46_66 11.551961
Rsp45_67 sp45_67 sp46_67 11.551961
Rsn45_67 sn45_67 sn46_67 11.551961
Rsp45_68 sp45_68 sp46_68 11.551961
Rsn45_68 sn45_68 sn46_68 11.551961
Rsp45_69 sp45_69 sp46_69 11.551961
Rsn45_69 sn45_69 sn46_69 11.551961
Rsp45_70 sp45_70 sp46_70 11.551961
Rsn45_70 sn45_70 sn46_70 11.551961
Rsp45_71 sp45_71 sp46_71 11.551961
Rsn45_71 sn45_71 sn46_71 11.551961
Rsp45_72 sp45_72 sp46_72 11.551961
Rsn45_72 sn45_72 sn46_72 11.551961
Rsp45_73 sp45_73 sp46_73 11.551961
Rsn45_73 sn45_73 sn46_73 11.551961
Rsp45_74 sp45_74 sp46_74 11.551961
Rsn45_74 sn45_74 sn46_74 11.551961
Rsp45_75 sp45_75 sp46_75 11.551961
Rsn45_75 sn45_75 sn46_75 11.551961
Rsp45_76 sp45_76 sp46_76 11.551961
Rsn45_76 sn45_76 sn46_76 11.551961
Rsp45_77 sp45_77 sp46_77 11.551961
Rsn45_77 sn45_77 sn46_77 11.551961
Rsp45_78 sp45_78 sp46_78 11.551961
Rsn45_78 sn45_78 sn46_78 11.551961
Rsp45_79 sp45_79 sp46_79 11.551961
Rsn45_79 sn45_79 sn46_79 11.551961
Rsp45_80 sp45_80 sp46_80 11.551961
Rsn45_80 sn45_80 sn46_80 11.551961
Rsp45_81 sp45_81 sp46_81 11.551961
Rsn45_81 sn45_81 sn46_81 11.551961
Rsp45_82 sp45_82 sp46_82 11.551961
Rsn45_82 sn45_82 sn46_82 11.551961
Rsp45_83 sp45_83 sp46_83 11.551961
Rsn45_83 sn45_83 sn46_83 11.551961
Rsp45_84 sp45_84 sp46_84 11.551961
Rsn45_84 sn45_84 sn46_84 11.551961
Rsp46_1 sp46_1 sp47_1 11.551961
Rsn46_1 sn46_1 sn47_1 11.551961
Rsp46_2 sp46_2 sp47_2 11.551961
Rsn46_2 sn46_2 sn47_2 11.551961
Rsp46_3 sp46_3 sp47_3 11.551961
Rsn46_3 sn46_3 sn47_3 11.551961
Rsp46_4 sp46_4 sp47_4 11.551961
Rsn46_4 sn46_4 sn47_4 11.551961
Rsp46_5 sp46_5 sp47_5 11.551961
Rsn46_5 sn46_5 sn47_5 11.551961
Rsp46_6 sp46_6 sp47_6 11.551961
Rsn46_6 sn46_6 sn47_6 11.551961
Rsp46_7 sp46_7 sp47_7 11.551961
Rsn46_7 sn46_7 sn47_7 11.551961
Rsp46_8 sp46_8 sp47_8 11.551961
Rsn46_8 sn46_8 sn47_8 11.551961
Rsp46_9 sp46_9 sp47_9 11.551961
Rsn46_9 sn46_9 sn47_9 11.551961
Rsp46_10 sp46_10 sp47_10 11.551961
Rsn46_10 sn46_10 sn47_10 11.551961
Rsp46_11 sp46_11 sp47_11 11.551961
Rsn46_11 sn46_11 sn47_11 11.551961
Rsp46_12 sp46_12 sp47_12 11.551961
Rsn46_12 sn46_12 sn47_12 11.551961
Rsp46_13 sp46_13 sp47_13 11.551961
Rsn46_13 sn46_13 sn47_13 11.551961
Rsp46_14 sp46_14 sp47_14 11.551961
Rsn46_14 sn46_14 sn47_14 11.551961
Rsp46_15 sp46_15 sp47_15 11.551961
Rsn46_15 sn46_15 sn47_15 11.551961
Rsp46_16 sp46_16 sp47_16 11.551961
Rsn46_16 sn46_16 sn47_16 11.551961
Rsp46_17 sp46_17 sp47_17 11.551961
Rsn46_17 sn46_17 sn47_17 11.551961
Rsp46_18 sp46_18 sp47_18 11.551961
Rsn46_18 sn46_18 sn47_18 11.551961
Rsp46_19 sp46_19 sp47_19 11.551961
Rsn46_19 sn46_19 sn47_19 11.551961
Rsp46_20 sp46_20 sp47_20 11.551961
Rsn46_20 sn46_20 sn47_20 11.551961
Rsp46_21 sp46_21 sp47_21 11.551961
Rsn46_21 sn46_21 sn47_21 11.551961
Rsp46_22 sp46_22 sp47_22 11.551961
Rsn46_22 sn46_22 sn47_22 11.551961
Rsp46_23 sp46_23 sp47_23 11.551961
Rsn46_23 sn46_23 sn47_23 11.551961
Rsp46_24 sp46_24 sp47_24 11.551961
Rsn46_24 sn46_24 sn47_24 11.551961
Rsp46_25 sp46_25 sp47_25 11.551961
Rsn46_25 sn46_25 sn47_25 11.551961
Rsp46_26 sp46_26 sp47_26 11.551961
Rsn46_26 sn46_26 sn47_26 11.551961
Rsp46_27 sp46_27 sp47_27 11.551961
Rsn46_27 sn46_27 sn47_27 11.551961
Rsp46_28 sp46_28 sp47_28 11.551961
Rsn46_28 sn46_28 sn47_28 11.551961
Rsp46_29 sp46_29 sp47_29 11.551961
Rsn46_29 sn46_29 sn47_29 11.551961
Rsp46_30 sp46_30 sp47_30 11.551961
Rsn46_30 sn46_30 sn47_30 11.551961
Rsp46_31 sp46_31 sp47_31 11.551961
Rsn46_31 sn46_31 sn47_31 11.551961
Rsp46_32 sp46_32 sp47_32 11.551961
Rsn46_32 sn46_32 sn47_32 11.551961
Rsp46_33 sp46_33 sp47_33 11.551961
Rsn46_33 sn46_33 sn47_33 11.551961
Rsp46_34 sp46_34 sp47_34 11.551961
Rsn46_34 sn46_34 sn47_34 11.551961
Rsp46_35 sp46_35 sp47_35 11.551961
Rsn46_35 sn46_35 sn47_35 11.551961
Rsp46_36 sp46_36 sp47_36 11.551961
Rsn46_36 sn46_36 sn47_36 11.551961
Rsp46_37 sp46_37 sp47_37 11.551961
Rsn46_37 sn46_37 sn47_37 11.551961
Rsp46_38 sp46_38 sp47_38 11.551961
Rsn46_38 sn46_38 sn47_38 11.551961
Rsp46_39 sp46_39 sp47_39 11.551961
Rsn46_39 sn46_39 sn47_39 11.551961
Rsp46_40 sp46_40 sp47_40 11.551961
Rsn46_40 sn46_40 sn47_40 11.551961
Rsp46_41 sp46_41 sp47_41 11.551961
Rsn46_41 sn46_41 sn47_41 11.551961
Rsp46_42 sp46_42 sp47_42 11.551961
Rsn46_42 sn46_42 sn47_42 11.551961
Rsp46_43 sp46_43 sp47_43 11.551961
Rsn46_43 sn46_43 sn47_43 11.551961
Rsp46_44 sp46_44 sp47_44 11.551961
Rsn46_44 sn46_44 sn47_44 11.551961
Rsp46_45 sp46_45 sp47_45 11.551961
Rsn46_45 sn46_45 sn47_45 11.551961
Rsp46_46 sp46_46 sp47_46 11.551961
Rsn46_46 sn46_46 sn47_46 11.551961
Rsp46_47 sp46_47 sp47_47 11.551961
Rsn46_47 sn46_47 sn47_47 11.551961
Rsp46_48 sp46_48 sp47_48 11.551961
Rsn46_48 sn46_48 sn47_48 11.551961
Rsp46_49 sp46_49 sp47_49 11.551961
Rsn46_49 sn46_49 sn47_49 11.551961
Rsp46_50 sp46_50 sp47_50 11.551961
Rsn46_50 sn46_50 sn47_50 11.551961
Rsp46_51 sp46_51 sp47_51 11.551961
Rsn46_51 sn46_51 sn47_51 11.551961
Rsp46_52 sp46_52 sp47_52 11.551961
Rsn46_52 sn46_52 sn47_52 11.551961
Rsp46_53 sp46_53 sp47_53 11.551961
Rsn46_53 sn46_53 sn47_53 11.551961
Rsp46_54 sp46_54 sp47_54 11.551961
Rsn46_54 sn46_54 sn47_54 11.551961
Rsp46_55 sp46_55 sp47_55 11.551961
Rsn46_55 sn46_55 sn47_55 11.551961
Rsp46_56 sp46_56 sp47_56 11.551961
Rsn46_56 sn46_56 sn47_56 11.551961
Rsp46_57 sp46_57 sp47_57 11.551961
Rsn46_57 sn46_57 sn47_57 11.551961
Rsp46_58 sp46_58 sp47_58 11.551961
Rsn46_58 sn46_58 sn47_58 11.551961
Rsp46_59 sp46_59 sp47_59 11.551961
Rsn46_59 sn46_59 sn47_59 11.551961
Rsp46_60 sp46_60 sp47_60 11.551961
Rsn46_60 sn46_60 sn47_60 11.551961
Rsp46_61 sp46_61 sp47_61 11.551961
Rsn46_61 sn46_61 sn47_61 11.551961
Rsp46_62 sp46_62 sp47_62 11.551961
Rsn46_62 sn46_62 sn47_62 11.551961
Rsp46_63 sp46_63 sp47_63 11.551961
Rsn46_63 sn46_63 sn47_63 11.551961
Rsp46_64 sp46_64 sp47_64 11.551961
Rsn46_64 sn46_64 sn47_64 11.551961
Rsp46_65 sp46_65 sp47_65 11.551961
Rsn46_65 sn46_65 sn47_65 11.551961
Rsp46_66 sp46_66 sp47_66 11.551961
Rsn46_66 sn46_66 sn47_66 11.551961
Rsp46_67 sp46_67 sp47_67 11.551961
Rsn46_67 sn46_67 sn47_67 11.551961
Rsp46_68 sp46_68 sp47_68 11.551961
Rsn46_68 sn46_68 sn47_68 11.551961
Rsp46_69 sp46_69 sp47_69 11.551961
Rsn46_69 sn46_69 sn47_69 11.551961
Rsp46_70 sp46_70 sp47_70 11.551961
Rsn46_70 sn46_70 sn47_70 11.551961
Rsp46_71 sp46_71 sp47_71 11.551961
Rsn46_71 sn46_71 sn47_71 11.551961
Rsp46_72 sp46_72 sp47_72 11.551961
Rsn46_72 sn46_72 sn47_72 11.551961
Rsp46_73 sp46_73 sp47_73 11.551961
Rsn46_73 sn46_73 sn47_73 11.551961
Rsp46_74 sp46_74 sp47_74 11.551961
Rsn46_74 sn46_74 sn47_74 11.551961
Rsp46_75 sp46_75 sp47_75 11.551961
Rsn46_75 sn46_75 sn47_75 11.551961
Rsp46_76 sp46_76 sp47_76 11.551961
Rsn46_76 sn46_76 sn47_76 11.551961
Rsp46_77 sp46_77 sp47_77 11.551961
Rsn46_77 sn46_77 sn47_77 11.551961
Rsp46_78 sp46_78 sp47_78 11.551961
Rsn46_78 sn46_78 sn47_78 11.551961
Rsp46_79 sp46_79 sp47_79 11.551961
Rsn46_79 sn46_79 sn47_79 11.551961
Rsp46_80 sp46_80 sp47_80 11.551961
Rsn46_80 sn46_80 sn47_80 11.551961
Rsp46_81 sp46_81 sp47_81 11.551961
Rsn46_81 sn46_81 sn47_81 11.551961
Rsp46_82 sp46_82 sp47_82 11.551961
Rsn46_82 sn46_82 sn47_82 11.551961
Rsp46_83 sp46_83 sp47_83 11.551961
Rsn46_83 sn46_83 sn47_83 11.551961
Rsp46_84 sp46_84 sp47_84 11.551961
Rsn46_84 sn46_84 sn47_84 11.551961
Rsp47_1 sp47_1 sp48_1 11.551961
Rsn47_1 sn47_1 sn48_1 11.551961
Rsp47_2 sp47_2 sp48_2 11.551961
Rsn47_2 sn47_2 sn48_2 11.551961
Rsp47_3 sp47_3 sp48_3 11.551961
Rsn47_3 sn47_3 sn48_3 11.551961
Rsp47_4 sp47_4 sp48_4 11.551961
Rsn47_4 sn47_4 sn48_4 11.551961
Rsp47_5 sp47_5 sp48_5 11.551961
Rsn47_5 sn47_5 sn48_5 11.551961
Rsp47_6 sp47_6 sp48_6 11.551961
Rsn47_6 sn47_6 sn48_6 11.551961
Rsp47_7 sp47_7 sp48_7 11.551961
Rsn47_7 sn47_7 sn48_7 11.551961
Rsp47_8 sp47_8 sp48_8 11.551961
Rsn47_8 sn47_8 sn48_8 11.551961
Rsp47_9 sp47_9 sp48_9 11.551961
Rsn47_9 sn47_9 sn48_9 11.551961
Rsp47_10 sp47_10 sp48_10 11.551961
Rsn47_10 sn47_10 sn48_10 11.551961
Rsp47_11 sp47_11 sp48_11 11.551961
Rsn47_11 sn47_11 sn48_11 11.551961
Rsp47_12 sp47_12 sp48_12 11.551961
Rsn47_12 sn47_12 sn48_12 11.551961
Rsp47_13 sp47_13 sp48_13 11.551961
Rsn47_13 sn47_13 sn48_13 11.551961
Rsp47_14 sp47_14 sp48_14 11.551961
Rsn47_14 sn47_14 sn48_14 11.551961
Rsp47_15 sp47_15 sp48_15 11.551961
Rsn47_15 sn47_15 sn48_15 11.551961
Rsp47_16 sp47_16 sp48_16 11.551961
Rsn47_16 sn47_16 sn48_16 11.551961
Rsp47_17 sp47_17 sp48_17 11.551961
Rsn47_17 sn47_17 sn48_17 11.551961
Rsp47_18 sp47_18 sp48_18 11.551961
Rsn47_18 sn47_18 sn48_18 11.551961
Rsp47_19 sp47_19 sp48_19 11.551961
Rsn47_19 sn47_19 sn48_19 11.551961
Rsp47_20 sp47_20 sp48_20 11.551961
Rsn47_20 sn47_20 sn48_20 11.551961
Rsp47_21 sp47_21 sp48_21 11.551961
Rsn47_21 sn47_21 sn48_21 11.551961
Rsp47_22 sp47_22 sp48_22 11.551961
Rsn47_22 sn47_22 sn48_22 11.551961
Rsp47_23 sp47_23 sp48_23 11.551961
Rsn47_23 sn47_23 sn48_23 11.551961
Rsp47_24 sp47_24 sp48_24 11.551961
Rsn47_24 sn47_24 sn48_24 11.551961
Rsp47_25 sp47_25 sp48_25 11.551961
Rsn47_25 sn47_25 sn48_25 11.551961
Rsp47_26 sp47_26 sp48_26 11.551961
Rsn47_26 sn47_26 sn48_26 11.551961
Rsp47_27 sp47_27 sp48_27 11.551961
Rsn47_27 sn47_27 sn48_27 11.551961
Rsp47_28 sp47_28 sp48_28 11.551961
Rsn47_28 sn47_28 sn48_28 11.551961
Rsp47_29 sp47_29 sp48_29 11.551961
Rsn47_29 sn47_29 sn48_29 11.551961
Rsp47_30 sp47_30 sp48_30 11.551961
Rsn47_30 sn47_30 sn48_30 11.551961
Rsp47_31 sp47_31 sp48_31 11.551961
Rsn47_31 sn47_31 sn48_31 11.551961
Rsp47_32 sp47_32 sp48_32 11.551961
Rsn47_32 sn47_32 sn48_32 11.551961
Rsp47_33 sp47_33 sp48_33 11.551961
Rsn47_33 sn47_33 sn48_33 11.551961
Rsp47_34 sp47_34 sp48_34 11.551961
Rsn47_34 sn47_34 sn48_34 11.551961
Rsp47_35 sp47_35 sp48_35 11.551961
Rsn47_35 sn47_35 sn48_35 11.551961
Rsp47_36 sp47_36 sp48_36 11.551961
Rsn47_36 sn47_36 sn48_36 11.551961
Rsp47_37 sp47_37 sp48_37 11.551961
Rsn47_37 sn47_37 sn48_37 11.551961
Rsp47_38 sp47_38 sp48_38 11.551961
Rsn47_38 sn47_38 sn48_38 11.551961
Rsp47_39 sp47_39 sp48_39 11.551961
Rsn47_39 sn47_39 sn48_39 11.551961
Rsp47_40 sp47_40 sp48_40 11.551961
Rsn47_40 sn47_40 sn48_40 11.551961
Rsp47_41 sp47_41 sp48_41 11.551961
Rsn47_41 sn47_41 sn48_41 11.551961
Rsp47_42 sp47_42 sp48_42 11.551961
Rsn47_42 sn47_42 sn48_42 11.551961
Rsp47_43 sp47_43 sp48_43 11.551961
Rsn47_43 sn47_43 sn48_43 11.551961
Rsp47_44 sp47_44 sp48_44 11.551961
Rsn47_44 sn47_44 sn48_44 11.551961
Rsp47_45 sp47_45 sp48_45 11.551961
Rsn47_45 sn47_45 sn48_45 11.551961
Rsp47_46 sp47_46 sp48_46 11.551961
Rsn47_46 sn47_46 sn48_46 11.551961
Rsp47_47 sp47_47 sp48_47 11.551961
Rsn47_47 sn47_47 sn48_47 11.551961
Rsp47_48 sp47_48 sp48_48 11.551961
Rsn47_48 sn47_48 sn48_48 11.551961
Rsp47_49 sp47_49 sp48_49 11.551961
Rsn47_49 sn47_49 sn48_49 11.551961
Rsp47_50 sp47_50 sp48_50 11.551961
Rsn47_50 sn47_50 sn48_50 11.551961
Rsp47_51 sp47_51 sp48_51 11.551961
Rsn47_51 sn47_51 sn48_51 11.551961
Rsp47_52 sp47_52 sp48_52 11.551961
Rsn47_52 sn47_52 sn48_52 11.551961
Rsp47_53 sp47_53 sp48_53 11.551961
Rsn47_53 sn47_53 sn48_53 11.551961
Rsp47_54 sp47_54 sp48_54 11.551961
Rsn47_54 sn47_54 sn48_54 11.551961
Rsp47_55 sp47_55 sp48_55 11.551961
Rsn47_55 sn47_55 sn48_55 11.551961
Rsp47_56 sp47_56 sp48_56 11.551961
Rsn47_56 sn47_56 sn48_56 11.551961
Rsp47_57 sp47_57 sp48_57 11.551961
Rsn47_57 sn47_57 sn48_57 11.551961
Rsp47_58 sp47_58 sp48_58 11.551961
Rsn47_58 sn47_58 sn48_58 11.551961
Rsp47_59 sp47_59 sp48_59 11.551961
Rsn47_59 sn47_59 sn48_59 11.551961
Rsp47_60 sp47_60 sp48_60 11.551961
Rsn47_60 sn47_60 sn48_60 11.551961
Rsp47_61 sp47_61 sp48_61 11.551961
Rsn47_61 sn47_61 sn48_61 11.551961
Rsp47_62 sp47_62 sp48_62 11.551961
Rsn47_62 sn47_62 sn48_62 11.551961
Rsp47_63 sp47_63 sp48_63 11.551961
Rsn47_63 sn47_63 sn48_63 11.551961
Rsp47_64 sp47_64 sp48_64 11.551961
Rsn47_64 sn47_64 sn48_64 11.551961
Rsp47_65 sp47_65 sp48_65 11.551961
Rsn47_65 sn47_65 sn48_65 11.551961
Rsp47_66 sp47_66 sp48_66 11.551961
Rsn47_66 sn47_66 sn48_66 11.551961
Rsp47_67 sp47_67 sp48_67 11.551961
Rsn47_67 sn47_67 sn48_67 11.551961
Rsp47_68 sp47_68 sp48_68 11.551961
Rsn47_68 sn47_68 sn48_68 11.551961
Rsp47_69 sp47_69 sp48_69 11.551961
Rsn47_69 sn47_69 sn48_69 11.551961
Rsp47_70 sp47_70 sp48_70 11.551961
Rsn47_70 sn47_70 sn48_70 11.551961
Rsp47_71 sp47_71 sp48_71 11.551961
Rsn47_71 sn47_71 sn48_71 11.551961
Rsp47_72 sp47_72 sp48_72 11.551961
Rsn47_72 sn47_72 sn48_72 11.551961
Rsp47_73 sp47_73 sp48_73 11.551961
Rsn47_73 sn47_73 sn48_73 11.551961
Rsp47_74 sp47_74 sp48_74 11.551961
Rsn47_74 sn47_74 sn48_74 11.551961
Rsp47_75 sp47_75 sp48_75 11.551961
Rsn47_75 sn47_75 sn48_75 11.551961
Rsp47_76 sp47_76 sp48_76 11.551961
Rsn47_76 sn47_76 sn48_76 11.551961
Rsp47_77 sp47_77 sp48_77 11.551961
Rsn47_77 sn47_77 sn48_77 11.551961
Rsp47_78 sp47_78 sp48_78 11.551961
Rsn47_78 sn47_78 sn48_78 11.551961
Rsp47_79 sp47_79 sp48_79 11.551961
Rsn47_79 sn47_79 sn48_79 11.551961
Rsp47_80 sp47_80 sp48_80 11.551961
Rsn47_80 sn47_80 sn48_80 11.551961
Rsp47_81 sp47_81 sp48_81 11.551961
Rsn47_81 sn47_81 sn48_81 11.551961
Rsp47_82 sp47_82 sp48_82 11.551961
Rsn47_82 sn47_82 sn48_82 11.551961
Rsp47_83 sp47_83 sp48_83 11.551961
Rsn47_83 sn47_83 sn48_83 11.551961
Rsp47_84 sp47_84 sp48_84 11.551961
Rsn47_84 sn47_84 sn48_84 11.551961
Rsp48_1 sp48_1 sp49_1 11.551961
Rsn48_1 sn48_1 sn49_1 11.551961
Rsp48_2 sp48_2 sp49_2 11.551961
Rsn48_2 sn48_2 sn49_2 11.551961
Rsp48_3 sp48_3 sp49_3 11.551961
Rsn48_3 sn48_3 sn49_3 11.551961
Rsp48_4 sp48_4 sp49_4 11.551961
Rsn48_4 sn48_4 sn49_4 11.551961
Rsp48_5 sp48_5 sp49_5 11.551961
Rsn48_5 sn48_5 sn49_5 11.551961
Rsp48_6 sp48_6 sp49_6 11.551961
Rsn48_6 sn48_6 sn49_6 11.551961
Rsp48_7 sp48_7 sp49_7 11.551961
Rsn48_7 sn48_7 sn49_7 11.551961
Rsp48_8 sp48_8 sp49_8 11.551961
Rsn48_8 sn48_8 sn49_8 11.551961
Rsp48_9 sp48_9 sp49_9 11.551961
Rsn48_9 sn48_9 sn49_9 11.551961
Rsp48_10 sp48_10 sp49_10 11.551961
Rsn48_10 sn48_10 sn49_10 11.551961
Rsp48_11 sp48_11 sp49_11 11.551961
Rsn48_11 sn48_11 sn49_11 11.551961
Rsp48_12 sp48_12 sp49_12 11.551961
Rsn48_12 sn48_12 sn49_12 11.551961
Rsp48_13 sp48_13 sp49_13 11.551961
Rsn48_13 sn48_13 sn49_13 11.551961
Rsp48_14 sp48_14 sp49_14 11.551961
Rsn48_14 sn48_14 sn49_14 11.551961
Rsp48_15 sp48_15 sp49_15 11.551961
Rsn48_15 sn48_15 sn49_15 11.551961
Rsp48_16 sp48_16 sp49_16 11.551961
Rsn48_16 sn48_16 sn49_16 11.551961
Rsp48_17 sp48_17 sp49_17 11.551961
Rsn48_17 sn48_17 sn49_17 11.551961
Rsp48_18 sp48_18 sp49_18 11.551961
Rsn48_18 sn48_18 sn49_18 11.551961
Rsp48_19 sp48_19 sp49_19 11.551961
Rsn48_19 sn48_19 sn49_19 11.551961
Rsp48_20 sp48_20 sp49_20 11.551961
Rsn48_20 sn48_20 sn49_20 11.551961
Rsp48_21 sp48_21 sp49_21 11.551961
Rsn48_21 sn48_21 sn49_21 11.551961
Rsp48_22 sp48_22 sp49_22 11.551961
Rsn48_22 sn48_22 sn49_22 11.551961
Rsp48_23 sp48_23 sp49_23 11.551961
Rsn48_23 sn48_23 sn49_23 11.551961
Rsp48_24 sp48_24 sp49_24 11.551961
Rsn48_24 sn48_24 sn49_24 11.551961
Rsp48_25 sp48_25 sp49_25 11.551961
Rsn48_25 sn48_25 sn49_25 11.551961
Rsp48_26 sp48_26 sp49_26 11.551961
Rsn48_26 sn48_26 sn49_26 11.551961
Rsp48_27 sp48_27 sp49_27 11.551961
Rsn48_27 sn48_27 sn49_27 11.551961
Rsp48_28 sp48_28 sp49_28 11.551961
Rsn48_28 sn48_28 sn49_28 11.551961
Rsp48_29 sp48_29 sp49_29 11.551961
Rsn48_29 sn48_29 sn49_29 11.551961
Rsp48_30 sp48_30 sp49_30 11.551961
Rsn48_30 sn48_30 sn49_30 11.551961
Rsp48_31 sp48_31 sp49_31 11.551961
Rsn48_31 sn48_31 sn49_31 11.551961
Rsp48_32 sp48_32 sp49_32 11.551961
Rsn48_32 sn48_32 sn49_32 11.551961
Rsp48_33 sp48_33 sp49_33 11.551961
Rsn48_33 sn48_33 sn49_33 11.551961
Rsp48_34 sp48_34 sp49_34 11.551961
Rsn48_34 sn48_34 sn49_34 11.551961
Rsp48_35 sp48_35 sp49_35 11.551961
Rsn48_35 sn48_35 sn49_35 11.551961
Rsp48_36 sp48_36 sp49_36 11.551961
Rsn48_36 sn48_36 sn49_36 11.551961
Rsp48_37 sp48_37 sp49_37 11.551961
Rsn48_37 sn48_37 sn49_37 11.551961
Rsp48_38 sp48_38 sp49_38 11.551961
Rsn48_38 sn48_38 sn49_38 11.551961
Rsp48_39 sp48_39 sp49_39 11.551961
Rsn48_39 sn48_39 sn49_39 11.551961
Rsp48_40 sp48_40 sp49_40 11.551961
Rsn48_40 sn48_40 sn49_40 11.551961
Rsp48_41 sp48_41 sp49_41 11.551961
Rsn48_41 sn48_41 sn49_41 11.551961
Rsp48_42 sp48_42 sp49_42 11.551961
Rsn48_42 sn48_42 sn49_42 11.551961
Rsp48_43 sp48_43 sp49_43 11.551961
Rsn48_43 sn48_43 sn49_43 11.551961
Rsp48_44 sp48_44 sp49_44 11.551961
Rsn48_44 sn48_44 sn49_44 11.551961
Rsp48_45 sp48_45 sp49_45 11.551961
Rsn48_45 sn48_45 sn49_45 11.551961
Rsp48_46 sp48_46 sp49_46 11.551961
Rsn48_46 sn48_46 sn49_46 11.551961
Rsp48_47 sp48_47 sp49_47 11.551961
Rsn48_47 sn48_47 sn49_47 11.551961
Rsp48_48 sp48_48 sp49_48 11.551961
Rsn48_48 sn48_48 sn49_48 11.551961
Rsp48_49 sp48_49 sp49_49 11.551961
Rsn48_49 sn48_49 sn49_49 11.551961
Rsp48_50 sp48_50 sp49_50 11.551961
Rsn48_50 sn48_50 sn49_50 11.551961
Rsp48_51 sp48_51 sp49_51 11.551961
Rsn48_51 sn48_51 sn49_51 11.551961
Rsp48_52 sp48_52 sp49_52 11.551961
Rsn48_52 sn48_52 sn49_52 11.551961
Rsp48_53 sp48_53 sp49_53 11.551961
Rsn48_53 sn48_53 sn49_53 11.551961
Rsp48_54 sp48_54 sp49_54 11.551961
Rsn48_54 sn48_54 sn49_54 11.551961
Rsp48_55 sp48_55 sp49_55 11.551961
Rsn48_55 sn48_55 sn49_55 11.551961
Rsp48_56 sp48_56 sp49_56 11.551961
Rsn48_56 sn48_56 sn49_56 11.551961
Rsp48_57 sp48_57 sp49_57 11.551961
Rsn48_57 sn48_57 sn49_57 11.551961
Rsp48_58 sp48_58 sp49_58 11.551961
Rsn48_58 sn48_58 sn49_58 11.551961
Rsp48_59 sp48_59 sp49_59 11.551961
Rsn48_59 sn48_59 sn49_59 11.551961
Rsp48_60 sp48_60 sp49_60 11.551961
Rsn48_60 sn48_60 sn49_60 11.551961
Rsp48_61 sp48_61 sp49_61 11.551961
Rsn48_61 sn48_61 sn49_61 11.551961
Rsp48_62 sp48_62 sp49_62 11.551961
Rsn48_62 sn48_62 sn49_62 11.551961
Rsp48_63 sp48_63 sp49_63 11.551961
Rsn48_63 sn48_63 sn49_63 11.551961
Rsp48_64 sp48_64 sp49_64 11.551961
Rsn48_64 sn48_64 sn49_64 11.551961
Rsp48_65 sp48_65 sp49_65 11.551961
Rsn48_65 sn48_65 sn49_65 11.551961
Rsp48_66 sp48_66 sp49_66 11.551961
Rsn48_66 sn48_66 sn49_66 11.551961
Rsp48_67 sp48_67 sp49_67 11.551961
Rsn48_67 sn48_67 sn49_67 11.551961
Rsp48_68 sp48_68 sp49_68 11.551961
Rsn48_68 sn48_68 sn49_68 11.551961
Rsp48_69 sp48_69 sp49_69 11.551961
Rsn48_69 sn48_69 sn49_69 11.551961
Rsp48_70 sp48_70 sp49_70 11.551961
Rsn48_70 sn48_70 sn49_70 11.551961
Rsp48_71 sp48_71 sp49_71 11.551961
Rsn48_71 sn48_71 sn49_71 11.551961
Rsp48_72 sp48_72 sp49_72 11.551961
Rsn48_72 sn48_72 sn49_72 11.551961
Rsp48_73 sp48_73 sp49_73 11.551961
Rsn48_73 sn48_73 sn49_73 11.551961
Rsp48_74 sp48_74 sp49_74 11.551961
Rsn48_74 sn48_74 sn49_74 11.551961
Rsp48_75 sp48_75 sp49_75 11.551961
Rsn48_75 sn48_75 sn49_75 11.551961
Rsp48_76 sp48_76 sp49_76 11.551961
Rsn48_76 sn48_76 sn49_76 11.551961
Rsp48_77 sp48_77 sp49_77 11.551961
Rsn48_77 sn48_77 sn49_77 11.551961
Rsp48_78 sp48_78 sp49_78 11.551961
Rsn48_78 sn48_78 sn49_78 11.551961
Rsp48_79 sp48_79 sp49_79 11.551961
Rsn48_79 sn48_79 sn49_79 11.551961
Rsp48_80 sp48_80 sp49_80 11.551961
Rsn48_80 sn48_80 sn49_80 11.551961
Rsp48_81 sp48_81 sp49_81 11.551961
Rsn48_81 sn48_81 sn49_81 11.551961
Rsp48_82 sp48_82 sp49_82 11.551961
Rsn48_82 sn48_82 sn49_82 11.551961
Rsp48_83 sp48_83 sp49_83 11.551961
Rsn48_83 sn48_83 sn49_83 11.551961
Rsp48_84 sp48_84 sp49_84 11.551961
Rsn48_84 sn48_84 sn49_84 11.551961
Rsp49_1 sp49_1 sp50_1 11.551961
Rsn49_1 sn49_1 sn50_1 11.551961
Rsp49_2 sp49_2 sp50_2 11.551961
Rsn49_2 sn49_2 sn50_2 11.551961
Rsp49_3 sp49_3 sp50_3 11.551961
Rsn49_3 sn49_3 sn50_3 11.551961
Rsp49_4 sp49_4 sp50_4 11.551961
Rsn49_4 sn49_4 sn50_4 11.551961
Rsp49_5 sp49_5 sp50_5 11.551961
Rsn49_5 sn49_5 sn50_5 11.551961
Rsp49_6 sp49_6 sp50_6 11.551961
Rsn49_6 sn49_6 sn50_6 11.551961
Rsp49_7 sp49_7 sp50_7 11.551961
Rsn49_7 sn49_7 sn50_7 11.551961
Rsp49_8 sp49_8 sp50_8 11.551961
Rsn49_8 sn49_8 sn50_8 11.551961
Rsp49_9 sp49_9 sp50_9 11.551961
Rsn49_9 sn49_9 sn50_9 11.551961
Rsp49_10 sp49_10 sp50_10 11.551961
Rsn49_10 sn49_10 sn50_10 11.551961
Rsp49_11 sp49_11 sp50_11 11.551961
Rsn49_11 sn49_11 sn50_11 11.551961
Rsp49_12 sp49_12 sp50_12 11.551961
Rsn49_12 sn49_12 sn50_12 11.551961
Rsp49_13 sp49_13 sp50_13 11.551961
Rsn49_13 sn49_13 sn50_13 11.551961
Rsp49_14 sp49_14 sp50_14 11.551961
Rsn49_14 sn49_14 sn50_14 11.551961
Rsp49_15 sp49_15 sp50_15 11.551961
Rsn49_15 sn49_15 sn50_15 11.551961
Rsp49_16 sp49_16 sp50_16 11.551961
Rsn49_16 sn49_16 sn50_16 11.551961
Rsp49_17 sp49_17 sp50_17 11.551961
Rsn49_17 sn49_17 sn50_17 11.551961
Rsp49_18 sp49_18 sp50_18 11.551961
Rsn49_18 sn49_18 sn50_18 11.551961
Rsp49_19 sp49_19 sp50_19 11.551961
Rsn49_19 sn49_19 sn50_19 11.551961
Rsp49_20 sp49_20 sp50_20 11.551961
Rsn49_20 sn49_20 sn50_20 11.551961
Rsp49_21 sp49_21 sp50_21 11.551961
Rsn49_21 sn49_21 sn50_21 11.551961
Rsp49_22 sp49_22 sp50_22 11.551961
Rsn49_22 sn49_22 sn50_22 11.551961
Rsp49_23 sp49_23 sp50_23 11.551961
Rsn49_23 sn49_23 sn50_23 11.551961
Rsp49_24 sp49_24 sp50_24 11.551961
Rsn49_24 sn49_24 sn50_24 11.551961
Rsp49_25 sp49_25 sp50_25 11.551961
Rsn49_25 sn49_25 sn50_25 11.551961
Rsp49_26 sp49_26 sp50_26 11.551961
Rsn49_26 sn49_26 sn50_26 11.551961
Rsp49_27 sp49_27 sp50_27 11.551961
Rsn49_27 sn49_27 sn50_27 11.551961
Rsp49_28 sp49_28 sp50_28 11.551961
Rsn49_28 sn49_28 sn50_28 11.551961
Rsp49_29 sp49_29 sp50_29 11.551961
Rsn49_29 sn49_29 sn50_29 11.551961
Rsp49_30 sp49_30 sp50_30 11.551961
Rsn49_30 sn49_30 sn50_30 11.551961
Rsp49_31 sp49_31 sp50_31 11.551961
Rsn49_31 sn49_31 sn50_31 11.551961
Rsp49_32 sp49_32 sp50_32 11.551961
Rsn49_32 sn49_32 sn50_32 11.551961
Rsp49_33 sp49_33 sp50_33 11.551961
Rsn49_33 sn49_33 sn50_33 11.551961
Rsp49_34 sp49_34 sp50_34 11.551961
Rsn49_34 sn49_34 sn50_34 11.551961
Rsp49_35 sp49_35 sp50_35 11.551961
Rsn49_35 sn49_35 sn50_35 11.551961
Rsp49_36 sp49_36 sp50_36 11.551961
Rsn49_36 sn49_36 sn50_36 11.551961
Rsp49_37 sp49_37 sp50_37 11.551961
Rsn49_37 sn49_37 sn50_37 11.551961
Rsp49_38 sp49_38 sp50_38 11.551961
Rsn49_38 sn49_38 sn50_38 11.551961
Rsp49_39 sp49_39 sp50_39 11.551961
Rsn49_39 sn49_39 sn50_39 11.551961
Rsp49_40 sp49_40 sp50_40 11.551961
Rsn49_40 sn49_40 sn50_40 11.551961
Rsp49_41 sp49_41 sp50_41 11.551961
Rsn49_41 sn49_41 sn50_41 11.551961
Rsp49_42 sp49_42 sp50_42 11.551961
Rsn49_42 sn49_42 sn50_42 11.551961
Rsp49_43 sp49_43 sp50_43 11.551961
Rsn49_43 sn49_43 sn50_43 11.551961
Rsp49_44 sp49_44 sp50_44 11.551961
Rsn49_44 sn49_44 sn50_44 11.551961
Rsp49_45 sp49_45 sp50_45 11.551961
Rsn49_45 sn49_45 sn50_45 11.551961
Rsp49_46 sp49_46 sp50_46 11.551961
Rsn49_46 sn49_46 sn50_46 11.551961
Rsp49_47 sp49_47 sp50_47 11.551961
Rsn49_47 sn49_47 sn50_47 11.551961
Rsp49_48 sp49_48 sp50_48 11.551961
Rsn49_48 sn49_48 sn50_48 11.551961
Rsp49_49 sp49_49 sp50_49 11.551961
Rsn49_49 sn49_49 sn50_49 11.551961
Rsp49_50 sp49_50 sp50_50 11.551961
Rsn49_50 sn49_50 sn50_50 11.551961
Rsp49_51 sp49_51 sp50_51 11.551961
Rsn49_51 sn49_51 sn50_51 11.551961
Rsp49_52 sp49_52 sp50_52 11.551961
Rsn49_52 sn49_52 sn50_52 11.551961
Rsp49_53 sp49_53 sp50_53 11.551961
Rsn49_53 sn49_53 sn50_53 11.551961
Rsp49_54 sp49_54 sp50_54 11.551961
Rsn49_54 sn49_54 sn50_54 11.551961
Rsp49_55 sp49_55 sp50_55 11.551961
Rsn49_55 sn49_55 sn50_55 11.551961
Rsp49_56 sp49_56 sp50_56 11.551961
Rsn49_56 sn49_56 sn50_56 11.551961
Rsp49_57 sp49_57 sp50_57 11.551961
Rsn49_57 sn49_57 sn50_57 11.551961
Rsp49_58 sp49_58 sp50_58 11.551961
Rsn49_58 sn49_58 sn50_58 11.551961
Rsp49_59 sp49_59 sp50_59 11.551961
Rsn49_59 sn49_59 sn50_59 11.551961
Rsp49_60 sp49_60 sp50_60 11.551961
Rsn49_60 sn49_60 sn50_60 11.551961
Rsp49_61 sp49_61 sp50_61 11.551961
Rsn49_61 sn49_61 sn50_61 11.551961
Rsp49_62 sp49_62 sp50_62 11.551961
Rsn49_62 sn49_62 sn50_62 11.551961
Rsp49_63 sp49_63 sp50_63 11.551961
Rsn49_63 sn49_63 sn50_63 11.551961
Rsp49_64 sp49_64 sp50_64 11.551961
Rsn49_64 sn49_64 sn50_64 11.551961
Rsp49_65 sp49_65 sp50_65 11.551961
Rsn49_65 sn49_65 sn50_65 11.551961
Rsp49_66 sp49_66 sp50_66 11.551961
Rsn49_66 sn49_66 sn50_66 11.551961
Rsp49_67 sp49_67 sp50_67 11.551961
Rsn49_67 sn49_67 sn50_67 11.551961
Rsp49_68 sp49_68 sp50_68 11.551961
Rsn49_68 sn49_68 sn50_68 11.551961
Rsp49_69 sp49_69 sp50_69 11.551961
Rsn49_69 sn49_69 sn50_69 11.551961
Rsp49_70 sp49_70 sp50_70 11.551961
Rsn49_70 sn49_70 sn50_70 11.551961
Rsp49_71 sp49_71 sp50_71 11.551961
Rsn49_71 sn49_71 sn50_71 11.551961
Rsp49_72 sp49_72 sp50_72 11.551961
Rsn49_72 sn49_72 sn50_72 11.551961
Rsp49_73 sp49_73 sp50_73 11.551961
Rsn49_73 sn49_73 sn50_73 11.551961
Rsp49_74 sp49_74 sp50_74 11.551961
Rsn49_74 sn49_74 sn50_74 11.551961
Rsp49_75 sp49_75 sp50_75 11.551961
Rsn49_75 sn49_75 sn50_75 11.551961
Rsp49_76 sp49_76 sp50_76 11.551961
Rsn49_76 sn49_76 sn50_76 11.551961
Rsp49_77 sp49_77 sp50_77 11.551961
Rsn49_77 sn49_77 sn50_77 11.551961
Rsp49_78 sp49_78 sp50_78 11.551961
Rsn49_78 sn49_78 sn50_78 11.551961
Rsp49_79 sp49_79 sp50_79 11.551961
Rsn49_79 sn49_79 sn50_79 11.551961
Rsp49_80 sp49_80 sp50_80 11.551961
Rsn49_80 sn49_80 sn50_80 11.551961
Rsp49_81 sp49_81 sp50_81 11.551961
Rsn49_81 sn49_81 sn50_81 11.551961
Rsp49_82 sp49_82 sp50_82 11.551961
Rsn49_82 sn49_82 sn50_82 11.551961
Rsp49_83 sp49_83 sp50_83 11.551961
Rsn49_83 sn49_83 sn50_83 11.551961
Rsp49_84 sp49_84 sp50_84 11.551961
Rsn49_84 sn49_84 sn50_84 11.551961
Rsp50_1 sp50_1 sp51_1 11.551961
Rsn50_1 sn50_1 sn51_1 11.551961
Rsp50_2 sp50_2 sp51_2 11.551961
Rsn50_2 sn50_2 sn51_2 11.551961
Rsp50_3 sp50_3 sp51_3 11.551961
Rsn50_3 sn50_3 sn51_3 11.551961
Rsp50_4 sp50_4 sp51_4 11.551961
Rsn50_4 sn50_4 sn51_4 11.551961
Rsp50_5 sp50_5 sp51_5 11.551961
Rsn50_5 sn50_5 sn51_5 11.551961
Rsp50_6 sp50_6 sp51_6 11.551961
Rsn50_6 sn50_6 sn51_6 11.551961
Rsp50_7 sp50_7 sp51_7 11.551961
Rsn50_7 sn50_7 sn51_7 11.551961
Rsp50_8 sp50_8 sp51_8 11.551961
Rsn50_8 sn50_8 sn51_8 11.551961
Rsp50_9 sp50_9 sp51_9 11.551961
Rsn50_9 sn50_9 sn51_9 11.551961
Rsp50_10 sp50_10 sp51_10 11.551961
Rsn50_10 sn50_10 sn51_10 11.551961
Rsp50_11 sp50_11 sp51_11 11.551961
Rsn50_11 sn50_11 sn51_11 11.551961
Rsp50_12 sp50_12 sp51_12 11.551961
Rsn50_12 sn50_12 sn51_12 11.551961
Rsp50_13 sp50_13 sp51_13 11.551961
Rsn50_13 sn50_13 sn51_13 11.551961
Rsp50_14 sp50_14 sp51_14 11.551961
Rsn50_14 sn50_14 sn51_14 11.551961
Rsp50_15 sp50_15 sp51_15 11.551961
Rsn50_15 sn50_15 sn51_15 11.551961
Rsp50_16 sp50_16 sp51_16 11.551961
Rsn50_16 sn50_16 sn51_16 11.551961
Rsp50_17 sp50_17 sp51_17 11.551961
Rsn50_17 sn50_17 sn51_17 11.551961
Rsp50_18 sp50_18 sp51_18 11.551961
Rsn50_18 sn50_18 sn51_18 11.551961
Rsp50_19 sp50_19 sp51_19 11.551961
Rsn50_19 sn50_19 sn51_19 11.551961
Rsp50_20 sp50_20 sp51_20 11.551961
Rsn50_20 sn50_20 sn51_20 11.551961
Rsp50_21 sp50_21 sp51_21 11.551961
Rsn50_21 sn50_21 sn51_21 11.551961
Rsp50_22 sp50_22 sp51_22 11.551961
Rsn50_22 sn50_22 sn51_22 11.551961
Rsp50_23 sp50_23 sp51_23 11.551961
Rsn50_23 sn50_23 sn51_23 11.551961
Rsp50_24 sp50_24 sp51_24 11.551961
Rsn50_24 sn50_24 sn51_24 11.551961
Rsp50_25 sp50_25 sp51_25 11.551961
Rsn50_25 sn50_25 sn51_25 11.551961
Rsp50_26 sp50_26 sp51_26 11.551961
Rsn50_26 sn50_26 sn51_26 11.551961
Rsp50_27 sp50_27 sp51_27 11.551961
Rsn50_27 sn50_27 sn51_27 11.551961
Rsp50_28 sp50_28 sp51_28 11.551961
Rsn50_28 sn50_28 sn51_28 11.551961
Rsp50_29 sp50_29 sp51_29 11.551961
Rsn50_29 sn50_29 sn51_29 11.551961
Rsp50_30 sp50_30 sp51_30 11.551961
Rsn50_30 sn50_30 sn51_30 11.551961
Rsp50_31 sp50_31 sp51_31 11.551961
Rsn50_31 sn50_31 sn51_31 11.551961
Rsp50_32 sp50_32 sp51_32 11.551961
Rsn50_32 sn50_32 sn51_32 11.551961
Rsp50_33 sp50_33 sp51_33 11.551961
Rsn50_33 sn50_33 sn51_33 11.551961
Rsp50_34 sp50_34 sp51_34 11.551961
Rsn50_34 sn50_34 sn51_34 11.551961
Rsp50_35 sp50_35 sp51_35 11.551961
Rsn50_35 sn50_35 sn51_35 11.551961
Rsp50_36 sp50_36 sp51_36 11.551961
Rsn50_36 sn50_36 sn51_36 11.551961
Rsp50_37 sp50_37 sp51_37 11.551961
Rsn50_37 sn50_37 sn51_37 11.551961
Rsp50_38 sp50_38 sp51_38 11.551961
Rsn50_38 sn50_38 sn51_38 11.551961
Rsp50_39 sp50_39 sp51_39 11.551961
Rsn50_39 sn50_39 sn51_39 11.551961
Rsp50_40 sp50_40 sp51_40 11.551961
Rsn50_40 sn50_40 sn51_40 11.551961
Rsp50_41 sp50_41 sp51_41 11.551961
Rsn50_41 sn50_41 sn51_41 11.551961
Rsp50_42 sp50_42 sp51_42 11.551961
Rsn50_42 sn50_42 sn51_42 11.551961
Rsp50_43 sp50_43 sp51_43 11.551961
Rsn50_43 sn50_43 sn51_43 11.551961
Rsp50_44 sp50_44 sp51_44 11.551961
Rsn50_44 sn50_44 sn51_44 11.551961
Rsp50_45 sp50_45 sp51_45 11.551961
Rsn50_45 sn50_45 sn51_45 11.551961
Rsp50_46 sp50_46 sp51_46 11.551961
Rsn50_46 sn50_46 sn51_46 11.551961
Rsp50_47 sp50_47 sp51_47 11.551961
Rsn50_47 sn50_47 sn51_47 11.551961
Rsp50_48 sp50_48 sp51_48 11.551961
Rsn50_48 sn50_48 sn51_48 11.551961
Rsp50_49 sp50_49 sp51_49 11.551961
Rsn50_49 sn50_49 sn51_49 11.551961
Rsp50_50 sp50_50 sp51_50 11.551961
Rsn50_50 sn50_50 sn51_50 11.551961
Rsp50_51 sp50_51 sp51_51 11.551961
Rsn50_51 sn50_51 sn51_51 11.551961
Rsp50_52 sp50_52 sp51_52 11.551961
Rsn50_52 sn50_52 sn51_52 11.551961
Rsp50_53 sp50_53 sp51_53 11.551961
Rsn50_53 sn50_53 sn51_53 11.551961
Rsp50_54 sp50_54 sp51_54 11.551961
Rsn50_54 sn50_54 sn51_54 11.551961
Rsp50_55 sp50_55 sp51_55 11.551961
Rsn50_55 sn50_55 sn51_55 11.551961
Rsp50_56 sp50_56 sp51_56 11.551961
Rsn50_56 sn50_56 sn51_56 11.551961
Rsp50_57 sp50_57 sp51_57 11.551961
Rsn50_57 sn50_57 sn51_57 11.551961
Rsp50_58 sp50_58 sp51_58 11.551961
Rsn50_58 sn50_58 sn51_58 11.551961
Rsp50_59 sp50_59 sp51_59 11.551961
Rsn50_59 sn50_59 sn51_59 11.551961
Rsp50_60 sp50_60 sp51_60 11.551961
Rsn50_60 sn50_60 sn51_60 11.551961
Rsp50_61 sp50_61 sp51_61 11.551961
Rsn50_61 sn50_61 sn51_61 11.551961
Rsp50_62 sp50_62 sp51_62 11.551961
Rsn50_62 sn50_62 sn51_62 11.551961
Rsp50_63 sp50_63 sp51_63 11.551961
Rsn50_63 sn50_63 sn51_63 11.551961
Rsp50_64 sp50_64 sp51_64 11.551961
Rsn50_64 sn50_64 sn51_64 11.551961
Rsp50_65 sp50_65 sp51_65 11.551961
Rsn50_65 sn50_65 sn51_65 11.551961
Rsp50_66 sp50_66 sp51_66 11.551961
Rsn50_66 sn50_66 sn51_66 11.551961
Rsp50_67 sp50_67 sp51_67 11.551961
Rsn50_67 sn50_67 sn51_67 11.551961
Rsp50_68 sp50_68 sp51_68 11.551961
Rsn50_68 sn50_68 sn51_68 11.551961
Rsp50_69 sp50_69 sp51_69 11.551961
Rsn50_69 sn50_69 sn51_69 11.551961
Rsp50_70 sp50_70 sp51_70 11.551961
Rsn50_70 sn50_70 sn51_70 11.551961
Rsp50_71 sp50_71 sp51_71 11.551961
Rsn50_71 sn50_71 sn51_71 11.551961
Rsp50_72 sp50_72 sp51_72 11.551961
Rsn50_72 sn50_72 sn51_72 11.551961
Rsp50_73 sp50_73 sp51_73 11.551961
Rsn50_73 sn50_73 sn51_73 11.551961
Rsp50_74 sp50_74 sp51_74 11.551961
Rsn50_74 sn50_74 sn51_74 11.551961
Rsp50_75 sp50_75 sp51_75 11.551961
Rsn50_75 sn50_75 sn51_75 11.551961
Rsp50_76 sp50_76 sp51_76 11.551961
Rsn50_76 sn50_76 sn51_76 11.551961
Rsp50_77 sp50_77 sp51_77 11.551961
Rsn50_77 sn50_77 sn51_77 11.551961
Rsp50_78 sp50_78 sp51_78 11.551961
Rsn50_78 sn50_78 sn51_78 11.551961
Rsp50_79 sp50_79 sp51_79 11.551961
Rsn50_79 sn50_79 sn51_79 11.551961
Rsp50_80 sp50_80 sp51_80 11.551961
Rsn50_80 sn50_80 sn51_80 11.551961
Rsp50_81 sp50_81 sp51_81 11.551961
Rsn50_81 sn50_81 sn51_81 11.551961
Rsp50_82 sp50_82 sp51_82 11.551961
Rsn50_82 sn50_82 sn51_82 11.551961
Rsp50_83 sp50_83 sp51_83 11.551961
Rsn50_83 sn50_83 sn51_83 11.551961
Rsp50_84 sp50_84 sp51_84 11.551961
Rsn50_84 sn50_84 sn51_84 11.551961
Rsp51_1 sp51_1 sp52_1 11.551961
Rsn51_1 sn51_1 sn52_1 11.551961
Rsp51_2 sp51_2 sp52_2 11.551961
Rsn51_2 sn51_2 sn52_2 11.551961
Rsp51_3 sp51_3 sp52_3 11.551961
Rsn51_3 sn51_3 sn52_3 11.551961
Rsp51_4 sp51_4 sp52_4 11.551961
Rsn51_4 sn51_4 sn52_4 11.551961
Rsp51_5 sp51_5 sp52_5 11.551961
Rsn51_5 sn51_5 sn52_5 11.551961
Rsp51_6 sp51_6 sp52_6 11.551961
Rsn51_6 sn51_6 sn52_6 11.551961
Rsp51_7 sp51_7 sp52_7 11.551961
Rsn51_7 sn51_7 sn52_7 11.551961
Rsp51_8 sp51_8 sp52_8 11.551961
Rsn51_8 sn51_8 sn52_8 11.551961
Rsp51_9 sp51_9 sp52_9 11.551961
Rsn51_9 sn51_9 sn52_9 11.551961
Rsp51_10 sp51_10 sp52_10 11.551961
Rsn51_10 sn51_10 sn52_10 11.551961
Rsp51_11 sp51_11 sp52_11 11.551961
Rsn51_11 sn51_11 sn52_11 11.551961
Rsp51_12 sp51_12 sp52_12 11.551961
Rsn51_12 sn51_12 sn52_12 11.551961
Rsp51_13 sp51_13 sp52_13 11.551961
Rsn51_13 sn51_13 sn52_13 11.551961
Rsp51_14 sp51_14 sp52_14 11.551961
Rsn51_14 sn51_14 sn52_14 11.551961
Rsp51_15 sp51_15 sp52_15 11.551961
Rsn51_15 sn51_15 sn52_15 11.551961
Rsp51_16 sp51_16 sp52_16 11.551961
Rsn51_16 sn51_16 sn52_16 11.551961
Rsp51_17 sp51_17 sp52_17 11.551961
Rsn51_17 sn51_17 sn52_17 11.551961
Rsp51_18 sp51_18 sp52_18 11.551961
Rsn51_18 sn51_18 sn52_18 11.551961
Rsp51_19 sp51_19 sp52_19 11.551961
Rsn51_19 sn51_19 sn52_19 11.551961
Rsp51_20 sp51_20 sp52_20 11.551961
Rsn51_20 sn51_20 sn52_20 11.551961
Rsp51_21 sp51_21 sp52_21 11.551961
Rsn51_21 sn51_21 sn52_21 11.551961
Rsp51_22 sp51_22 sp52_22 11.551961
Rsn51_22 sn51_22 sn52_22 11.551961
Rsp51_23 sp51_23 sp52_23 11.551961
Rsn51_23 sn51_23 sn52_23 11.551961
Rsp51_24 sp51_24 sp52_24 11.551961
Rsn51_24 sn51_24 sn52_24 11.551961
Rsp51_25 sp51_25 sp52_25 11.551961
Rsn51_25 sn51_25 sn52_25 11.551961
Rsp51_26 sp51_26 sp52_26 11.551961
Rsn51_26 sn51_26 sn52_26 11.551961
Rsp51_27 sp51_27 sp52_27 11.551961
Rsn51_27 sn51_27 sn52_27 11.551961
Rsp51_28 sp51_28 sp52_28 11.551961
Rsn51_28 sn51_28 sn52_28 11.551961
Rsp51_29 sp51_29 sp52_29 11.551961
Rsn51_29 sn51_29 sn52_29 11.551961
Rsp51_30 sp51_30 sp52_30 11.551961
Rsn51_30 sn51_30 sn52_30 11.551961
Rsp51_31 sp51_31 sp52_31 11.551961
Rsn51_31 sn51_31 sn52_31 11.551961
Rsp51_32 sp51_32 sp52_32 11.551961
Rsn51_32 sn51_32 sn52_32 11.551961
Rsp51_33 sp51_33 sp52_33 11.551961
Rsn51_33 sn51_33 sn52_33 11.551961
Rsp51_34 sp51_34 sp52_34 11.551961
Rsn51_34 sn51_34 sn52_34 11.551961
Rsp51_35 sp51_35 sp52_35 11.551961
Rsn51_35 sn51_35 sn52_35 11.551961
Rsp51_36 sp51_36 sp52_36 11.551961
Rsn51_36 sn51_36 sn52_36 11.551961
Rsp51_37 sp51_37 sp52_37 11.551961
Rsn51_37 sn51_37 sn52_37 11.551961
Rsp51_38 sp51_38 sp52_38 11.551961
Rsn51_38 sn51_38 sn52_38 11.551961
Rsp51_39 sp51_39 sp52_39 11.551961
Rsn51_39 sn51_39 sn52_39 11.551961
Rsp51_40 sp51_40 sp52_40 11.551961
Rsn51_40 sn51_40 sn52_40 11.551961
Rsp51_41 sp51_41 sp52_41 11.551961
Rsn51_41 sn51_41 sn52_41 11.551961
Rsp51_42 sp51_42 sp52_42 11.551961
Rsn51_42 sn51_42 sn52_42 11.551961
Rsp51_43 sp51_43 sp52_43 11.551961
Rsn51_43 sn51_43 sn52_43 11.551961
Rsp51_44 sp51_44 sp52_44 11.551961
Rsn51_44 sn51_44 sn52_44 11.551961
Rsp51_45 sp51_45 sp52_45 11.551961
Rsn51_45 sn51_45 sn52_45 11.551961
Rsp51_46 sp51_46 sp52_46 11.551961
Rsn51_46 sn51_46 sn52_46 11.551961
Rsp51_47 sp51_47 sp52_47 11.551961
Rsn51_47 sn51_47 sn52_47 11.551961
Rsp51_48 sp51_48 sp52_48 11.551961
Rsn51_48 sn51_48 sn52_48 11.551961
Rsp51_49 sp51_49 sp52_49 11.551961
Rsn51_49 sn51_49 sn52_49 11.551961
Rsp51_50 sp51_50 sp52_50 11.551961
Rsn51_50 sn51_50 sn52_50 11.551961
Rsp51_51 sp51_51 sp52_51 11.551961
Rsn51_51 sn51_51 sn52_51 11.551961
Rsp51_52 sp51_52 sp52_52 11.551961
Rsn51_52 sn51_52 sn52_52 11.551961
Rsp51_53 sp51_53 sp52_53 11.551961
Rsn51_53 sn51_53 sn52_53 11.551961
Rsp51_54 sp51_54 sp52_54 11.551961
Rsn51_54 sn51_54 sn52_54 11.551961
Rsp51_55 sp51_55 sp52_55 11.551961
Rsn51_55 sn51_55 sn52_55 11.551961
Rsp51_56 sp51_56 sp52_56 11.551961
Rsn51_56 sn51_56 sn52_56 11.551961
Rsp51_57 sp51_57 sp52_57 11.551961
Rsn51_57 sn51_57 sn52_57 11.551961
Rsp51_58 sp51_58 sp52_58 11.551961
Rsn51_58 sn51_58 sn52_58 11.551961
Rsp51_59 sp51_59 sp52_59 11.551961
Rsn51_59 sn51_59 sn52_59 11.551961
Rsp51_60 sp51_60 sp52_60 11.551961
Rsn51_60 sn51_60 sn52_60 11.551961
Rsp51_61 sp51_61 sp52_61 11.551961
Rsn51_61 sn51_61 sn52_61 11.551961
Rsp51_62 sp51_62 sp52_62 11.551961
Rsn51_62 sn51_62 sn52_62 11.551961
Rsp51_63 sp51_63 sp52_63 11.551961
Rsn51_63 sn51_63 sn52_63 11.551961
Rsp51_64 sp51_64 sp52_64 11.551961
Rsn51_64 sn51_64 sn52_64 11.551961
Rsp51_65 sp51_65 sp52_65 11.551961
Rsn51_65 sn51_65 sn52_65 11.551961
Rsp51_66 sp51_66 sp52_66 11.551961
Rsn51_66 sn51_66 sn52_66 11.551961
Rsp51_67 sp51_67 sp52_67 11.551961
Rsn51_67 sn51_67 sn52_67 11.551961
Rsp51_68 sp51_68 sp52_68 11.551961
Rsn51_68 sn51_68 sn52_68 11.551961
Rsp51_69 sp51_69 sp52_69 11.551961
Rsn51_69 sn51_69 sn52_69 11.551961
Rsp51_70 sp51_70 sp52_70 11.551961
Rsn51_70 sn51_70 sn52_70 11.551961
Rsp51_71 sp51_71 sp52_71 11.551961
Rsn51_71 sn51_71 sn52_71 11.551961
Rsp51_72 sp51_72 sp52_72 11.551961
Rsn51_72 sn51_72 sn52_72 11.551961
Rsp51_73 sp51_73 sp52_73 11.551961
Rsn51_73 sn51_73 sn52_73 11.551961
Rsp51_74 sp51_74 sp52_74 11.551961
Rsn51_74 sn51_74 sn52_74 11.551961
Rsp51_75 sp51_75 sp52_75 11.551961
Rsn51_75 sn51_75 sn52_75 11.551961
Rsp51_76 sp51_76 sp52_76 11.551961
Rsn51_76 sn51_76 sn52_76 11.551961
Rsp51_77 sp51_77 sp52_77 11.551961
Rsn51_77 sn51_77 sn52_77 11.551961
Rsp51_78 sp51_78 sp52_78 11.551961
Rsn51_78 sn51_78 sn52_78 11.551961
Rsp51_79 sp51_79 sp52_79 11.551961
Rsn51_79 sn51_79 sn52_79 11.551961
Rsp51_80 sp51_80 sp52_80 11.551961
Rsn51_80 sn51_80 sn52_80 11.551961
Rsp51_81 sp51_81 sp52_81 11.551961
Rsn51_81 sn51_81 sn52_81 11.551961
Rsp51_82 sp51_82 sp52_82 11.551961
Rsn51_82 sn51_82 sn52_82 11.551961
Rsp51_83 sp51_83 sp52_83 11.551961
Rsn51_83 sn51_83 sn52_83 11.551961
Rsp51_84 sp51_84 sp52_84 11.551961
Rsn51_84 sn51_84 sn52_84 11.551961
Rsp52_1 sp52_1 sp53_1 11.551961
Rsn52_1 sn52_1 sn53_1 11.551961
Rsp52_2 sp52_2 sp53_2 11.551961
Rsn52_2 sn52_2 sn53_2 11.551961
Rsp52_3 sp52_3 sp53_3 11.551961
Rsn52_3 sn52_3 sn53_3 11.551961
Rsp52_4 sp52_4 sp53_4 11.551961
Rsn52_4 sn52_4 sn53_4 11.551961
Rsp52_5 sp52_5 sp53_5 11.551961
Rsn52_5 sn52_5 sn53_5 11.551961
Rsp52_6 sp52_6 sp53_6 11.551961
Rsn52_6 sn52_6 sn53_6 11.551961
Rsp52_7 sp52_7 sp53_7 11.551961
Rsn52_7 sn52_7 sn53_7 11.551961
Rsp52_8 sp52_8 sp53_8 11.551961
Rsn52_8 sn52_8 sn53_8 11.551961
Rsp52_9 sp52_9 sp53_9 11.551961
Rsn52_9 sn52_9 sn53_9 11.551961
Rsp52_10 sp52_10 sp53_10 11.551961
Rsn52_10 sn52_10 sn53_10 11.551961
Rsp52_11 sp52_11 sp53_11 11.551961
Rsn52_11 sn52_11 sn53_11 11.551961
Rsp52_12 sp52_12 sp53_12 11.551961
Rsn52_12 sn52_12 sn53_12 11.551961
Rsp52_13 sp52_13 sp53_13 11.551961
Rsn52_13 sn52_13 sn53_13 11.551961
Rsp52_14 sp52_14 sp53_14 11.551961
Rsn52_14 sn52_14 sn53_14 11.551961
Rsp52_15 sp52_15 sp53_15 11.551961
Rsn52_15 sn52_15 sn53_15 11.551961
Rsp52_16 sp52_16 sp53_16 11.551961
Rsn52_16 sn52_16 sn53_16 11.551961
Rsp52_17 sp52_17 sp53_17 11.551961
Rsn52_17 sn52_17 sn53_17 11.551961
Rsp52_18 sp52_18 sp53_18 11.551961
Rsn52_18 sn52_18 sn53_18 11.551961
Rsp52_19 sp52_19 sp53_19 11.551961
Rsn52_19 sn52_19 sn53_19 11.551961
Rsp52_20 sp52_20 sp53_20 11.551961
Rsn52_20 sn52_20 sn53_20 11.551961
Rsp52_21 sp52_21 sp53_21 11.551961
Rsn52_21 sn52_21 sn53_21 11.551961
Rsp52_22 sp52_22 sp53_22 11.551961
Rsn52_22 sn52_22 sn53_22 11.551961
Rsp52_23 sp52_23 sp53_23 11.551961
Rsn52_23 sn52_23 sn53_23 11.551961
Rsp52_24 sp52_24 sp53_24 11.551961
Rsn52_24 sn52_24 sn53_24 11.551961
Rsp52_25 sp52_25 sp53_25 11.551961
Rsn52_25 sn52_25 sn53_25 11.551961
Rsp52_26 sp52_26 sp53_26 11.551961
Rsn52_26 sn52_26 sn53_26 11.551961
Rsp52_27 sp52_27 sp53_27 11.551961
Rsn52_27 sn52_27 sn53_27 11.551961
Rsp52_28 sp52_28 sp53_28 11.551961
Rsn52_28 sn52_28 sn53_28 11.551961
Rsp52_29 sp52_29 sp53_29 11.551961
Rsn52_29 sn52_29 sn53_29 11.551961
Rsp52_30 sp52_30 sp53_30 11.551961
Rsn52_30 sn52_30 sn53_30 11.551961
Rsp52_31 sp52_31 sp53_31 11.551961
Rsn52_31 sn52_31 sn53_31 11.551961
Rsp52_32 sp52_32 sp53_32 11.551961
Rsn52_32 sn52_32 sn53_32 11.551961
Rsp52_33 sp52_33 sp53_33 11.551961
Rsn52_33 sn52_33 sn53_33 11.551961
Rsp52_34 sp52_34 sp53_34 11.551961
Rsn52_34 sn52_34 sn53_34 11.551961
Rsp52_35 sp52_35 sp53_35 11.551961
Rsn52_35 sn52_35 sn53_35 11.551961
Rsp52_36 sp52_36 sp53_36 11.551961
Rsn52_36 sn52_36 sn53_36 11.551961
Rsp52_37 sp52_37 sp53_37 11.551961
Rsn52_37 sn52_37 sn53_37 11.551961
Rsp52_38 sp52_38 sp53_38 11.551961
Rsn52_38 sn52_38 sn53_38 11.551961
Rsp52_39 sp52_39 sp53_39 11.551961
Rsn52_39 sn52_39 sn53_39 11.551961
Rsp52_40 sp52_40 sp53_40 11.551961
Rsn52_40 sn52_40 sn53_40 11.551961
Rsp52_41 sp52_41 sp53_41 11.551961
Rsn52_41 sn52_41 sn53_41 11.551961
Rsp52_42 sp52_42 sp53_42 11.551961
Rsn52_42 sn52_42 sn53_42 11.551961
Rsp52_43 sp52_43 sp53_43 11.551961
Rsn52_43 sn52_43 sn53_43 11.551961
Rsp52_44 sp52_44 sp53_44 11.551961
Rsn52_44 sn52_44 sn53_44 11.551961
Rsp52_45 sp52_45 sp53_45 11.551961
Rsn52_45 sn52_45 sn53_45 11.551961
Rsp52_46 sp52_46 sp53_46 11.551961
Rsn52_46 sn52_46 sn53_46 11.551961
Rsp52_47 sp52_47 sp53_47 11.551961
Rsn52_47 sn52_47 sn53_47 11.551961
Rsp52_48 sp52_48 sp53_48 11.551961
Rsn52_48 sn52_48 sn53_48 11.551961
Rsp52_49 sp52_49 sp53_49 11.551961
Rsn52_49 sn52_49 sn53_49 11.551961
Rsp52_50 sp52_50 sp53_50 11.551961
Rsn52_50 sn52_50 sn53_50 11.551961
Rsp52_51 sp52_51 sp53_51 11.551961
Rsn52_51 sn52_51 sn53_51 11.551961
Rsp52_52 sp52_52 sp53_52 11.551961
Rsn52_52 sn52_52 sn53_52 11.551961
Rsp52_53 sp52_53 sp53_53 11.551961
Rsn52_53 sn52_53 sn53_53 11.551961
Rsp52_54 sp52_54 sp53_54 11.551961
Rsn52_54 sn52_54 sn53_54 11.551961
Rsp52_55 sp52_55 sp53_55 11.551961
Rsn52_55 sn52_55 sn53_55 11.551961
Rsp52_56 sp52_56 sp53_56 11.551961
Rsn52_56 sn52_56 sn53_56 11.551961
Rsp52_57 sp52_57 sp53_57 11.551961
Rsn52_57 sn52_57 sn53_57 11.551961
Rsp52_58 sp52_58 sp53_58 11.551961
Rsn52_58 sn52_58 sn53_58 11.551961
Rsp52_59 sp52_59 sp53_59 11.551961
Rsn52_59 sn52_59 sn53_59 11.551961
Rsp52_60 sp52_60 sp53_60 11.551961
Rsn52_60 sn52_60 sn53_60 11.551961
Rsp52_61 sp52_61 sp53_61 11.551961
Rsn52_61 sn52_61 sn53_61 11.551961
Rsp52_62 sp52_62 sp53_62 11.551961
Rsn52_62 sn52_62 sn53_62 11.551961
Rsp52_63 sp52_63 sp53_63 11.551961
Rsn52_63 sn52_63 sn53_63 11.551961
Rsp52_64 sp52_64 sp53_64 11.551961
Rsn52_64 sn52_64 sn53_64 11.551961
Rsp52_65 sp52_65 sp53_65 11.551961
Rsn52_65 sn52_65 sn53_65 11.551961
Rsp52_66 sp52_66 sp53_66 11.551961
Rsn52_66 sn52_66 sn53_66 11.551961
Rsp52_67 sp52_67 sp53_67 11.551961
Rsn52_67 sn52_67 sn53_67 11.551961
Rsp52_68 sp52_68 sp53_68 11.551961
Rsn52_68 sn52_68 sn53_68 11.551961
Rsp52_69 sp52_69 sp53_69 11.551961
Rsn52_69 sn52_69 sn53_69 11.551961
Rsp52_70 sp52_70 sp53_70 11.551961
Rsn52_70 sn52_70 sn53_70 11.551961
Rsp52_71 sp52_71 sp53_71 11.551961
Rsn52_71 sn52_71 sn53_71 11.551961
Rsp52_72 sp52_72 sp53_72 11.551961
Rsn52_72 sn52_72 sn53_72 11.551961
Rsp52_73 sp52_73 sp53_73 11.551961
Rsn52_73 sn52_73 sn53_73 11.551961
Rsp52_74 sp52_74 sp53_74 11.551961
Rsn52_74 sn52_74 sn53_74 11.551961
Rsp52_75 sp52_75 sp53_75 11.551961
Rsn52_75 sn52_75 sn53_75 11.551961
Rsp52_76 sp52_76 sp53_76 11.551961
Rsn52_76 sn52_76 sn53_76 11.551961
Rsp52_77 sp52_77 sp53_77 11.551961
Rsn52_77 sn52_77 sn53_77 11.551961
Rsp52_78 sp52_78 sp53_78 11.551961
Rsn52_78 sn52_78 sn53_78 11.551961
Rsp52_79 sp52_79 sp53_79 11.551961
Rsn52_79 sn52_79 sn53_79 11.551961
Rsp52_80 sp52_80 sp53_80 11.551961
Rsn52_80 sn52_80 sn53_80 11.551961
Rsp52_81 sp52_81 sp53_81 11.551961
Rsn52_81 sn52_81 sn53_81 11.551961
Rsp52_82 sp52_82 sp53_82 11.551961
Rsn52_82 sn52_82 sn53_82 11.551961
Rsp52_83 sp52_83 sp53_83 11.551961
Rsn52_83 sn52_83 sn53_83 11.551961
Rsp52_84 sp52_84 sp53_84 11.551961
Rsn52_84 sn52_84 sn53_84 11.551961
Rsp53_1 sp53_1 sp54_1 11.551961
Rsn53_1 sn53_1 sn54_1 11.551961
Rsp53_2 sp53_2 sp54_2 11.551961
Rsn53_2 sn53_2 sn54_2 11.551961
Rsp53_3 sp53_3 sp54_3 11.551961
Rsn53_3 sn53_3 sn54_3 11.551961
Rsp53_4 sp53_4 sp54_4 11.551961
Rsn53_4 sn53_4 sn54_4 11.551961
Rsp53_5 sp53_5 sp54_5 11.551961
Rsn53_5 sn53_5 sn54_5 11.551961
Rsp53_6 sp53_6 sp54_6 11.551961
Rsn53_6 sn53_6 sn54_6 11.551961
Rsp53_7 sp53_7 sp54_7 11.551961
Rsn53_7 sn53_7 sn54_7 11.551961
Rsp53_8 sp53_8 sp54_8 11.551961
Rsn53_8 sn53_8 sn54_8 11.551961
Rsp53_9 sp53_9 sp54_9 11.551961
Rsn53_9 sn53_9 sn54_9 11.551961
Rsp53_10 sp53_10 sp54_10 11.551961
Rsn53_10 sn53_10 sn54_10 11.551961
Rsp53_11 sp53_11 sp54_11 11.551961
Rsn53_11 sn53_11 sn54_11 11.551961
Rsp53_12 sp53_12 sp54_12 11.551961
Rsn53_12 sn53_12 sn54_12 11.551961
Rsp53_13 sp53_13 sp54_13 11.551961
Rsn53_13 sn53_13 sn54_13 11.551961
Rsp53_14 sp53_14 sp54_14 11.551961
Rsn53_14 sn53_14 sn54_14 11.551961
Rsp53_15 sp53_15 sp54_15 11.551961
Rsn53_15 sn53_15 sn54_15 11.551961
Rsp53_16 sp53_16 sp54_16 11.551961
Rsn53_16 sn53_16 sn54_16 11.551961
Rsp53_17 sp53_17 sp54_17 11.551961
Rsn53_17 sn53_17 sn54_17 11.551961
Rsp53_18 sp53_18 sp54_18 11.551961
Rsn53_18 sn53_18 sn54_18 11.551961
Rsp53_19 sp53_19 sp54_19 11.551961
Rsn53_19 sn53_19 sn54_19 11.551961
Rsp53_20 sp53_20 sp54_20 11.551961
Rsn53_20 sn53_20 sn54_20 11.551961
Rsp53_21 sp53_21 sp54_21 11.551961
Rsn53_21 sn53_21 sn54_21 11.551961
Rsp53_22 sp53_22 sp54_22 11.551961
Rsn53_22 sn53_22 sn54_22 11.551961
Rsp53_23 sp53_23 sp54_23 11.551961
Rsn53_23 sn53_23 sn54_23 11.551961
Rsp53_24 sp53_24 sp54_24 11.551961
Rsn53_24 sn53_24 sn54_24 11.551961
Rsp53_25 sp53_25 sp54_25 11.551961
Rsn53_25 sn53_25 sn54_25 11.551961
Rsp53_26 sp53_26 sp54_26 11.551961
Rsn53_26 sn53_26 sn54_26 11.551961
Rsp53_27 sp53_27 sp54_27 11.551961
Rsn53_27 sn53_27 sn54_27 11.551961
Rsp53_28 sp53_28 sp54_28 11.551961
Rsn53_28 sn53_28 sn54_28 11.551961
Rsp53_29 sp53_29 sp54_29 11.551961
Rsn53_29 sn53_29 sn54_29 11.551961
Rsp53_30 sp53_30 sp54_30 11.551961
Rsn53_30 sn53_30 sn54_30 11.551961
Rsp53_31 sp53_31 sp54_31 11.551961
Rsn53_31 sn53_31 sn54_31 11.551961
Rsp53_32 sp53_32 sp54_32 11.551961
Rsn53_32 sn53_32 sn54_32 11.551961
Rsp53_33 sp53_33 sp54_33 11.551961
Rsn53_33 sn53_33 sn54_33 11.551961
Rsp53_34 sp53_34 sp54_34 11.551961
Rsn53_34 sn53_34 sn54_34 11.551961
Rsp53_35 sp53_35 sp54_35 11.551961
Rsn53_35 sn53_35 sn54_35 11.551961
Rsp53_36 sp53_36 sp54_36 11.551961
Rsn53_36 sn53_36 sn54_36 11.551961
Rsp53_37 sp53_37 sp54_37 11.551961
Rsn53_37 sn53_37 sn54_37 11.551961
Rsp53_38 sp53_38 sp54_38 11.551961
Rsn53_38 sn53_38 sn54_38 11.551961
Rsp53_39 sp53_39 sp54_39 11.551961
Rsn53_39 sn53_39 sn54_39 11.551961
Rsp53_40 sp53_40 sp54_40 11.551961
Rsn53_40 sn53_40 sn54_40 11.551961
Rsp53_41 sp53_41 sp54_41 11.551961
Rsn53_41 sn53_41 sn54_41 11.551961
Rsp53_42 sp53_42 sp54_42 11.551961
Rsn53_42 sn53_42 sn54_42 11.551961
Rsp53_43 sp53_43 sp54_43 11.551961
Rsn53_43 sn53_43 sn54_43 11.551961
Rsp53_44 sp53_44 sp54_44 11.551961
Rsn53_44 sn53_44 sn54_44 11.551961
Rsp53_45 sp53_45 sp54_45 11.551961
Rsn53_45 sn53_45 sn54_45 11.551961
Rsp53_46 sp53_46 sp54_46 11.551961
Rsn53_46 sn53_46 sn54_46 11.551961
Rsp53_47 sp53_47 sp54_47 11.551961
Rsn53_47 sn53_47 sn54_47 11.551961
Rsp53_48 sp53_48 sp54_48 11.551961
Rsn53_48 sn53_48 sn54_48 11.551961
Rsp53_49 sp53_49 sp54_49 11.551961
Rsn53_49 sn53_49 sn54_49 11.551961
Rsp53_50 sp53_50 sp54_50 11.551961
Rsn53_50 sn53_50 sn54_50 11.551961
Rsp53_51 sp53_51 sp54_51 11.551961
Rsn53_51 sn53_51 sn54_51 11.551961
Rsp53_52 sp53_52 sp54_52 11.551961
Rsn53_52 sn53_52 sn54_52 11.551961
Rsp53_53 sp53_53 sp54_53 11.551961
Rsn53_53 sn53_53 sn54_53 11.551961
Rsp53_54 sp53_54 sp54_54 11.551961
Rsn53_54 sn53_54 sn54_54 11.551961
Rsp53_55 sp53_55 sp54_55 11.551961
Rsn53_55 sn53_55 sn54_55 11.551961
Rsp53_56 sp53_56 sp54_56 11.551961
Rsn53_56 sn53_56 sn54_56 11.551961
Rsp53_57 sp53_57 sp54_57 11.551961
Rsn53_57 sn53_57 sn54_57 11.551961
Rsp53_58 sp53_58 sp54_58 11.551961
Rsn53_58 sn53_58 sn54_58 11.551961
Rsp53_59 sp53_59 sp54_59 11.551961
Rsn53_59 sn53_59 sn54_59 11.551961
Rsp53_60 sp53_60 sp54_60 11.551961
Rsn53_60 sn53_60 sn54_60 11.551961
Rsp53_61 sp53_61 sp54_61 11.551961
Rsn53_61 sn53_61 sn54_61 11.551961
Rsp53_62 sp53_62 sp54_62 11.551961
Rsn53_62 sn53_62 sn54_62 11.551961
Rsp53_63 sp53_63 sp54_63 11.551961
Rsn53_63 sn53_63 sn54_63 11.551961
Rsp53_64 sp53_64 sp54_64 11.551961
Rsn53_64 sn53_64 sn54_64 11.551961
Rsp53_65 sp53_65 sp54_65 11.551961
Rsn53_65 sn53_65 sn54_65 11.551961
Rsp53_66 sp53_66 sp54_66 11.551961
Rsn53_66 sn53_66 sn54_66 11.551961
Rsp53_67 sp53_67 sp54_67 11.551961
Rsn53_67 sn53_67 sn54_67 11.551961
Rsp53_68 sp53_68 sp54_68 11.551961
Rsn53_68 sn53_68 sn54_68 11.551961
Rsp53_69 sp53_69 sp54_69 11.551961
Rsn53_69 sn53_69 sn54_69 11.551961
Rsp53_70 sp53_70 sp54_70 11.551961
Rsn53_70 sn53_70 sn54_70 11.551961
Rsp53_71 sp53_71 sp54_71 11.551961
Rsn53_71 sn53_71 sn54_71 11.551961
Rsp53_72 sp53_72 sp54_72 11.551961
Rsn53_72 sn53_72 sn54_72 11.551961
Rsp53_73 sp53_73 sp54_73 11.551961
Rsn53_73 sn53_73 sn54_73 11.551961
Rsp53_74 sp53_74 sp54_74 11.551961
Rsn53_74 sn53_74 sn54_74 11.551961
Rsp53_75 sp53_75 sp54_75 11.551961
Rsn53_75 sn53_75 sn54_75 11.551961
Rsp53_76 sp53_76 sp54_76 11.551961
Rsn53_76 sn53_76 sn54_76 11.551961
Rsp53_77 sp53_77 sp54_77 11.551961
Rsn53_77 sn53_77 sn54_77 11.551961
Rsp53_78 sp53_78 sp54_78 11.551961
Rsn53_78 sn53_78 sn54_78 11.551961
Rsp53_79 sp53_79 sp54_79 11.551961
Rsn53_79 sn53_79 sn54_79 11.551961
Rsp53_80 sp53_80 sp54_80 11.551961
Rsn53_80 sn53_80 sn54_80 11.551961
Rsp53_81 sp53_81 sp54_81 11.551961
Rsn53_81 sn53_81 sn54_81 11.551961
Rsp53_82 sp53_82 sp54_82 11.551961
Rsn53_82 sn53_82 sn54_82 11.551961
Rsp53_83 sp53_83 sp54_83 11.551961
Rsn53_83 sn53_83 sn54_83 11.551961
Rsp53_84 sp53_84 sp54_84 11.551961
Rsn53_84 sn53_84 sn54_84 11.551961
Rsp54_1 sp54_1 sp55_1 11.551961
Rsn54_1 sn54_1 sn55_1 11.551961
Rsp54_2 sp54_2 sp55_2 11.551961
Rsn54_2 sn54_2 sn55_2 11.551961
Rsp54_3 sp54_3 sp55_3 11.551961
Rsn54_3 sn54_3 sn55_3 11.551961
Rsp54_4 sp54_4 sp55_4 11.551961
Rsn54_4 sn54_4 sn55_4 11.551961
Rsp54_5 sp54_5 sp55_5 11.551961
Rsn54_5 sn54_5 sn55_5 11.551961
Rsp54_6 sp54_6 sp55_6 11.551961
Rsn54_6 sn54_6 sn55_6 11.551961
Rsp54_7 sp54_7 sp55_7 11.551961
Rsn54_7 sn54_7 sn55_7 11.551961
Rsp54_8 sp54_8 sp55_8 11.551961
Rsn54_8 sn54_8 sn55_8 11.551961
Rsp54_9 sp54_9 sp55_9 11.551961
Rsn54_9 sn54_9 sn55_9 11.551961
Rsp54_10 sp54_10 sp55_10 11.551961
Rsn54_10 sn54_10 sn55_10 11.551961
Rsp54_11 sp54_11 sp55_11 11.551961
Rsn54_11 sn54_11 sn55_11 11.551961
Rsp54_12 sp54_12 sp55_12 11.551961
Rsn54_12 sn54_12 sn55_12 11.551961
Rsp54_13 sp54_13 sp55_13 11.551961
Rsn54_13 sn54_13 sn55_13 11.551961
Rsp54_14 sp54_14 sp55_14 11.551961
Rsn54_14 sn54_14 sn55_14 11.551961
Rsp54_15 sp54_15 sp55_15 11.551961
Rsn54_15 sn54_15 sn55_15 11.551961
Rsp54_16 sp54_16 sp55_16 11.551961
Rsn54_16 sn54_16 sn55_16 11.551961
Rsp54_17 sp54_17 sp55_17 11.551961
Rsn54_17 sn54_17 sn55_17 11.551961
Rsp54_18 sp54_18 sp55_18 11.551961
Rsn54_18 sn54_18 sn55_18 11.551961
Rsp54_19 sp54_19 sp55_19 11.551961
Rsn54_19 sn54_19 sn55_19 11.551961
Rsp54_20 sp54_20 sp55_20 11.551961
Rsn54_20 sn54_20 sn55_20 11.551961
Rsp54_21 sp54_21 sp55_21 11.551961
Rsn54_21 sn54_21 sn55_21 11.551961
Rsp54_22 sp54_22 sp55_22 11.551961
Rsn54_22 sn54_22 sn55_22 11.551961
Rsp54_23 sp54_23 sp55_23 11.551961
Rsn54_23 sn54_23 sn55_23 11.551961
Rsp54_24 sp54_24 sp55_24 11.551961
Rsn54_24 sn54_24 sn55_24 11.551961
Rsp54_25 sp54_25 sp55_25 11.551961
Rsn54_25 sn54_25 sn55_25 11.551961
Rsp54_26 sp54_26 sp55_26 11.551961
Rsn54_26 sn54_26 sn55_26 11.551961
Rsp54_27 sp54_27 sp55_27 11.551961
Rsn54_27 sn54_27 sn55_27 11.551961
Rsp54_28 sp54_28 sp55_28 11.551961
Rsn54_28 sn54_28 sn55_28 11.551961
Rsp54_29 sp54_29 sp55_29 11.551961
Rsn54_29 sn54_29 sn55_29 11.551961
Rsp54_30 sp54_30 sp55_30 11.551961
Rsn54_30 sn54_30 sn55_30 11.551961
Rsp54_31 sp54_31 sp55_31 11.551961
Rsn54_31 sn54_31 sn55_31 11.551961
Rsp54_32 sp54_32 sp55_32 11.551961
Rsn54_32 sn54_32 sn55_32 11.551961
Rsp54_33 sp54_33 sp55_33 11.551961
Rsn54_33 sn54_33 sn55_33 11.551961
Rsp54_34 sp54_34 sp55_34 11.551961
Rsn54_34 sn54_34 sn55_34 11.551961
Rsp54_35 sp54_35 sp55_35 11.551961
Rsn54_35 sn54_35 sn55_35 11.551961
Rsp54_36 sp54_36 sp55_36 11.551961
Rsn54_36 sn54_36 sn55_36 11.551961
Rsp54_37 sp54_37 sp55_37 11.551961
Rsn54_37 sn54_37 sn55_37 11.551961
Rsp54_38 sp54_38 sp55_38 11.551961
Rsn54_38 sn54_38 sn55_38 11.551961
Rsp54_39 sp54_39 sp55_39 11.551961
Rsn54_39 sn54_39 sn55_39 11.551961
Rsp54_40 sp54_40 sp55_40 11.551961
Rsn54_40 sn54_40 sn55_40 11.551961
Rsp54_41 sp54_41 sp55_41 11.551961
Rsn54_41 sn54_41 sn55_41 11.551961
Rsp54_42 sp54_42 sp55_42 11.551961
Rsn54_42 sn54_42 sn55_42 11.551961
Rsp54_43 sp54_43 sp55_43 11.551961
Rsn54_43 sn54_43 sn55_43 11.551961
Rsp54_44 sp54_44 sp55_44 11.551961
Rsn54_44 sn54_44 sn55_44 11.551961
Rsp54_45 sp54_45 sp55_45 11.551961
Rsn54_45 sn54_45 sn55_45 11.551961
Rsp54_46 sp54_46 sp55_46 11.551961
Rsn54_46 sn54_46 sn55_46 11.551961
Rsp54_47 sp54_47 sp55_47 11.551961
Rsn54_47 sn54_47 sn55_47 11.551961
Rsp54_48 sp54_48 sp55_48 11.551961
Rsn54_48 sn54_48 sn55_48 11.551961
Rsp54_49 sp54_49 sp55_49 11.551961
Rsn54_49 sn54_49 sn55_49 11.551961
Rsp54_50 sp54_50 sp55_50 11.551961
Rsn54_50 sn54_50 sn55_50 11.551961
Rsp54_51 sp54_51 sp55_51 11.551961
Rsn54_51 sn54_51 sn55_51 11.551961
Rsp54_52 sp54_52 sp55_52 11.551961
Rsn54_52 sn54_52 sn55_52 11.551961
Rsp54_53 sp54_53 sp55_53 11.551961
Rsn54_53 sn54_53 sn55_53 11.551961
Rsp54_54 sp54_54 sp55_54 11.551961
Rsn54_54 sn54_54 sn55_54 11.551961
Rsp54_55 sp54_55 sp55_55 11.551961
Rsn54_55 sn54_55 sn55_55 11.551961
Rsp54_56 sp54_56 sp55_56 11.551961
Rsn54_56 sn54_56 sn55_56 11.551961
Rsp54_57 sp54_57 sp55_57 11.551961
Rsn54_57 sn54_57 sn55_57 11.551961
Rsp54_58 sp54_58 sp55_58 11.551961
Rsn54_58 sn54_58 sn55_58 11.551961
Rsp54_59 sp54_59 sp55_59 11.551961
Rsn54_59 sn54_59 sn55_59 11.551961
Rsp54_60 sp54_60 sp55_60 11.551961
Rsn54_60 sn54_60 sn55_60 11.551961
Rsp54_61 sp54_61 sp55_61 11.551961
Rsn54_61 sn54_61 sn55_61 11.551961
Rsp54_62 sp54_62 sp55_62 11.551961
Rsn54_62 sn54_62 sn55_62 11.551961
Rsp54_63 sp54_63 sp55_63 11.551961
Rsn54_63 sn54_63 sn55_63 11.551961
Rsp54_64 sp54_64 sp55_64 11.551961
Rsn54_64 sn54_64 sn55_64 11.551961
Rsp54_65 sp54_65 sp55_65 11.551961
Rsn54_65 sn54_65 sn55_65 11.551961
Rsp54_66 sp54_66 sp55_66 11.551961
Rsn54_66 sn54_66 sn55_66 11.551961
Rsp54_67 sp54_67 sp55_67 11.551961
Rsn54_67 sn54_67 sn55_67 11.551961
Rsp54_68 sp54_68 sp55_68 11.551961
Rsn54_68 sn54_68 sn55_68 11.551961
Rsp54_69 sp54_69 sp55_69 11.551961
Rsn54_69 sn54_69 sn55_69 11.551961
Rsp54_70 sp54_70 sp55_70 11.551961
Rsn54_70 sn54_70 sn55_70 11.551961
Rsp54_71 sp54_71 sp55_71 11.551961
Rsn54_71 sn54_71 sn55_71 11.551961
Rsp54_72 sp54_72 sp55_72 11.551961
Rsn54_72 sn54_72 sn55_72 11.551961
Rsp54_73 sp54_73 sp55_73 11.551961
Rsn54_73 sn54_73 sn55_73 11.551961
Rsp54_74 sp54_74 sp55_74 11.551961
Rsn54_74 sn54_74 sn55_74 11.551961
Rsp54_75 sp54_75 sp55_75 11.551961
Rsn54_75 sn54_75 sn55_75 11.551961
Rsp54_76 sp54_76 sp55_76 11.551961
Rsn54_76 sn54_76 sn55_76 11.551961
Rsp54_77 sp54_77 sp55_77 11.551961
Rsn54_77 sn54_77 sn55_77 11.551961
Rsp54_78 sp54_78 sp55_78 11.551961
Rsn54_78 sn54_78 sn55_78 11.551961
Rsp54_79 sp54_79 sp55_79 11.551961
Rsn54_79 sn54_79 sn55_79 11.551961
Rsp54_80 sp54_80 sp55_80 11.551961
Rsn54_80 sn54_80 sn55_80 11.551961
Rsp54_81 sp54_81 sp55_81 11.551961
Rsn54_81 sn54_81 sn55_81 11.551961
Rsp54_82 sp54_82 sp55_82 11.551961
Rsn54_82 sn54_82 sn55_82 11.551961
Rsp54_83 sp54_83 sp55_83 11.551961
Rsn54_83 sn54_83 sn55_83 11.551961
Rsp54_84 sp54_84 sp55_84 11.551961
Rsn54_84 sn54_84 sn55_84 11.551961
Rsp55_1 sp55_1 sp56_1 11.551961
Rsn55_1 sn55_1 sn56_1 11.551961
Rsp55_2 sp55_2 sp56_2 11.551961
Rsn55_2 sn55_2 sn56_2 11.551961
Rsp55_3 sp55_3 sp56_3 11.551961
Rsn55_3 sn55_3 sn56_3 11.551961
Rsp55_4 sp55_4 sp56_4 11.551961
Rsn55_4 sn55_4 sn56_4 11.551961
Rsp55_5 sp55_5 sp56_5 11.551961
Rsn55_5 sn55_5 sn56_5 11.551961
Rsp55_6 sp55_6 sp56_6 11.551961
Rsn55_6 sn55_6 sn56_6 11.551961
Rsp55_7 sp55_7 sp56_7 11.551961
Rsn55_7 sn55_7 sn56_7 11.551961
Rsp55_8 sp55_8 sp56_8 11.551961
Rsn55_8 sn55_8 sn56_8 11.551961
Rsp55_9 sp55_9 sp56_9 11.551961
Rsn55_9 sn55_9 sn56_9 11.551961
Rsp55_10 sp55_10 sp56_10 11.551961
Rsn55_10 sn55_10 sn56_10 11.551961
Rsp55_11 sp55_11 sp56_11 11.551961
Rsn55_11 sn55_11 sn56_11 11.551961
Rsp55_12 sp55_12 sp56_12 11.551961
Rsn55_12 sn55_12 sn56_12 11.551961
Rsp55_13 sp55_13 sp56_13 11.551961
Rsn55_13 sn55_13 sn56_13 11.551961
Rsp55_14 sp55_14 sp56_14 11.551961
Rsn55_14 sn55_14 sn56_14 11.551961
Rsp55_15 sp55_15 sp56_15 11.551961
Rsn55_15 sn55_15 sn56_15 11.551961
Rsp55_16 sp55_16 sp56_16 11.551961
Rsn55_16 sn55_16 sn56_16 11.551961
Rsp55_17 sp55_17 sp56_17 11.551961
Rsn55_17 sn55_17 sn56_17 11.551961
Rsp55_18 sp55_18 sp56_18 11.551961
Rsn55_18 sn55_18 sn56_18 11.551961
Rsp55_19 sp55_19 sp56_19 11.551961
Rsn55_19 sn55_19 sn56_19 11.551961
Rsp55_20 sp55_20 sp56_20 11.551961
Rsn55_20 sn55_20 sn56_20 11.551961
Rsp55_21 sp55_21 sp56_21 11.551961
Rsn55_21 sn55_21 sn56_21 11.551961
Rsp55_22 sp55_22 sp56_22 11.551961
Rsn55_22 sn55_22 sn56_22 11.551961
Rsp55_23 sp55_23 sp56_23 11.551961
Rsn55_23 sn55_23 sn56_23 11.551961
Rsp55_24 sp55_24 sp56_24 11.551961
Rsn55_24 sn55_24 sn56_24 11.551961
Rsp55_25 sp55_25 sp56_25 11.551961
Rsn55_25 sn55_25 sn56_25 11.551961
Rsp55_26 sp55_26 sp56_26 11.551961
Rsn55_26 sn55_26 sn56_26 11.551961
Rsp55_27 sp55_27 sp56_27 11.551961
Rsn55_27 sn55_27 sn56_27 11.551961
Rsp55_28 sp55_28 sp56_28 11.551961
Rsn55_28 sn55_28 sn56_28 11.551961
Rsp55_29 sp55_29 sp56_29 11.551961
Rsn55_29 sn55_29 sn56_29 11.551961
Rsp55_30 sp55_30 sp56_30 11.551961
Rsn55_30 sn55_30 sn56_30 11.551961
Rsp55_31 sp55_31 sp56_31 11.551961
Rsn55_31 sn55_31 sn56_31 11.551961
Rsp55_32 sp55_32 sp56_32 11.551961
Rsn55_32 sn55_32 sn56_32 11.551961
Rsp55_33 sp55_33 sp56_33 11.551961
Rsn55_33 sn55_33 sn56_33 11.551961
Rsp55_34 sp55_34 sp56_34 11.551961
Rsn55_34 sn55_34 sn56_34 11.551961
Rsp55_35 sp55_35 sp56_35 11.551961
Rsn55_35 sn55_35 sn56_35 11.551961
Rsp55_36 sp55_36 sp56_36 11.551961
Rsn55_36 sn55_36 sn56_36 11.551961
Rsp55_37 sp55_37 sp56_37 11.551961
Rsn55_37 sn55_37 sn56_37 11.551961
Rsp55_38 sp55_38 sp56_38 11.551961
Rsn55_38 sn55_38 sn56_38 11.551961
Rsp55_39 sp55_39 sp56_39 11.551961
Rsn55_39 sn55_39 sn56_39 11.551961
Rsp55_40 sp55_40 sp56_40 11.551961
Rsn55_40 sn55_40 sn56_40 11.551961
Rsp55_41 sp55_41 sp56_41 11.551961
Rsn55_41 sn55_41 sn56_41 11.551961
Rsp55_42 sp55_42 sp56_42 11.551961
Rsn55_42 sn55_42 sn56_42 11.551961
Rsp55_43 sp55_43 sp56_43 11.551961
Rsn55_43 sn55_43 sn56_43 11.551961
Rsp55_44 sp55_44 sp56_44 11.551961
Rsn55_44 sn55_44 sn56_44 11.551961
Rsp55_45 sp55_45 sp56_45 11.551961
Rsn55_45 sn55_45 sn56_45 11.551961
Rsp55_46 sp55_46 sp56_46 11.551961
Rsn55_46 sn55_46 sn56_46 11.551961
Rsp55_47 sp55_47 sp56_47 11.551961
Rsn55_47 sn55_47 sn56_47 11.551961
Rsp55_48 sp55_48 sp56_48 11.551961
Rsn55_48 sn55_48 sn56_48 11.551961
Rsp55_49 sp55_49 sp56_49 11.551961
Rsn55_49 sn55_49 sn56_49 11.551961
Rsp55_50 sp55_50 sp56_50 11.551961
Rsn55_50 sn55_50 sn56_50 11.551961
Rsp55_51 sp55_51 sp56_51 11.551961
Rsn55_51 sn55_51 sn56_51 11.551961
Rsp55_52 sp55_52 sp56_52 11.551961
Rsn55_52 sn55_52 sn56_52 11.551961
Rsp55_53 sp55_53 sp56_53 11.551961
Rsn55_53 sn55_53 sn56_53 11.551961
Rsp55_54 sp55_54 sp56_54 11.551961
Rsn55_54 sn55_54 sn56_54 11.551961
Rsp55_55 sp55_55 sp56_55 11.551961
Rsn55_55 sn55_55 sn56_55 11.551961
Rsp55_56 sp55_56 sp56_56 11.551961
Rsn55_56 sn55_56 sn56_56 11.551961
Rsp55_57 sp55_57 sp56_57 11.551961
Rsn55_57 sn55_57 sn56_57 11.551961
Rsp55_58 sp55_58 sp56_58 11.551961
Rsn55_58 sn55_58 sn56_58 11.551961
Rsp55_59 sp55_59 sp56_59 11.551961
Rsn55_59 sn55_59 sn56_59 11.551961
Rsp55_60 sp55_60 sp56_60 11.551961
Rsn55_60 sn55_60 sn56_60 11.551961
Rsp55_61 sp55_61 sp56_61 11.551961
Rsn55_61 sn55_61 sn56_61 11.551961
Rsp55_62 sp55_62 sp56_62 11.551961
Rsn55_62 sn55_62 sn56_62 11.551961
Rsp55_63 sp55_63 sp56_63 11.551961
Rsn55_63 sn55_63 sn56_63 11.551961
Rsp55_64 sp55_64 sp56_64 11.551961
Rsn55_64 sn55_64 sn56_64 11.551961
Rsp55_65 sp55_65 sp56_65 11.551961
Rsn55_65 sn55_65 sn56_65 11.551961
Rsp55_66 sp55_66 sp56_66 11.551961
Rsn55_66 sn55_66 sn56_66 11.551961
Rsp55_67 sp55_67 sp56_67 11.551961
Rsn55_67 sn55_67 sn56_67 11.551961
Rsp55_68 sp55_68 sp56_68 11.551961
Rsn55_68 sn55_68 sn56_68 11.551961
Rsp55_69 sp55_69 sp56_69 11.551961
Rsn55_69 sn55_69 sn56_69 11.551961
Rsp55_70 sp55_70 sp56_70 11.551961
Rsn55_70 sn55_70 sn56_70 11.551961
Rsp55_71 sp55_71 sp56_71 11.551961
Rsn55_71 sn55_71 sn56_71 11.551961
Rsp55_72 sp55_72 sp56_72 11.551961
Rsn55_72 sn55_72 sn56_72 11.551961
Rsp55_73 sp55_73 sp56_73 11.551961
Rsn55_73 sn55_73 sn56_73 11.551961
Rsp55_74 sp55_74 sp56_74 11.551961
Rsn55_74 sn55_74 sn56_74 11.551961
Rsp55_75 sp55_75 sp56_75 11.551961
Rsn55_75 sn55_75 sn56_75 11.551961
Rsp55_76 sp55_76 sp56_76 11.551961
Rsn55_76 sn55_76 sn56_76 11.551961
Rsp55_77 sp55_77 sp56_77 11.551961
Rsn55_77 sn55_77 sn56_77 11.551961
Rsp55_78 sp55_78 sp56_78 11.551961
Rsn55_78 sn55_78 sn56_78 11.551961
Rsp55_79 sp55_79 sp56_79 11.551961
Rsn55_79 sn55_79 sn56_79 11.551961
Rsp55_80 sp55_80 sp56_80 11.551961
Rsn55_80 sn55_80 sn56_80 11.551961
Rsp55_81 sp55_81 sp56_81 11.551961
Rsn55_81 sn55_81 sn56_81 11.551961
Rsp55_82 sp55_82 sp56_82 11.551961
Rsn55_82 sn55_82 sn56_82 11.551961
Rsp55_83 sp55_83 sp56_83 11.551961
Rsn55_83 sn55_83 sn56_83 11.551961
Rsp55_84 sp55_84 sp56_84 11.551961
Rsn55_84 sn55_84 sn56_84 11.551961
Rsp56_1 sp56_1 sp57_1 11.551961
Rsn56_1 sn56_1 sn57_1 11.551961
Rsp56_2 sp56_2 sp57_2 11.551961
Rsn56_2 sn56_2 sn57_2 11.551961
Rsp56_3 sp56_3 sp57_3 11.551961
Rsn56_3 sn56_3 sn57_3 11.551961
Rsp56_4 sp56_4 sp57_4 11.551961
Rsn56_4 sn56_4 sn57_4 11.551961
Rsp56_5 sp56_5 sp57_5 11.551961
Rsn56_5 sn56_5 sn57_5 11.551961
Rsp56_6 sp56_6 sp57_6 11.551961
Rsn56_6 sn56_6 sn57_6 11.551961
Rsp56_7 sp56_7 sp57_7 11.551961
Rsn56_7 sn56_7 sn57_7 11.551961
Rsp56_8 sp56_8 sp57_8 11.551961
Rsn56_8 sn56_8 sn57_8 11.551961
Rsp56_9 sp56_9 sp57_9 11.551961
Rsn56_9 sn56_9 sn57_9 11.551961
Rsp56_10 sp56_10 sp57_10 11.551961
Rsn56_10 sn56_10 sn57_10 11.551961
Rsp56_11 sp56_11 sp57_11 11.551961
Rsn56_11 sn56_11 sn57_11 11.551961
Rsp56_12 sp56_12 sp57_12 11.551961
Rsn56_12 sn56_12 sn57_12 11.551961
Rsp56_13 sp56_13 sp57_13 11.551961
Rsn56_13 sn56_13 sn57_13 11.551961
Rsp56_14 sp56_14 sp57_14 11.551961
Rsn56_14 sn56_14 sn57_14 11.551961
Rsp56_15 sp56_15 sp57_15 11.551961
Rsn56_15 sn56_15 sn57_15 11.551961
Rsp56_16 sp56_16 sp57_16 11.551961
Rsn56_16 sn56_16 sn57_16 11.551961
Rsp56_17 sp56_17 sp57_17 11.551961
Rsn56_17 sn56_17 sn57_17 11.551961
Rsp56_18 sp56_18 sp57_18 11.551961
Rsn56_18 sn56_18 sn57_18 11.551961
Rsp56_19 sp56_19 sp57_19 11.551961
Rsn56_19 sn56_19 sn57_19 11.551961
Rsp56_20 sp56_20 sp57_20 11.551961
Rsn56_20 sn56_20 sn57_20 11.551961
Rsp56_21 sp56_21 sp57_21 11.551961
Rsn56_21 sn56_21 sn57_21 11.551961
Rsp56_22 sp56_22 sp57_22 11.551961
Rsn56_22 sn56_22 sn57_22 11.551961
Rsp56_23 sp56_23 sp57_23 11.551961
Rsn56_23 sn56_23 sn57_23 11.551961
Rsp56_24 sp56_24 sp57_24 11.551961
Rsn56_24 sn56_24 sn57_24 11.551961
Rsp56_25 sp56_25 sp57_25 11.551961
Rsn56_25 sn56_25 sn57_25 11.551961
Rsp56_26 sp56_26 sp57_26 11.551961
Rsn56_26 sn56_26 sn57_26 11.551961
Rsp56_27 sp56_27 sp57_27 11.551961
Rsn56_27 sn56_27 sn57_27 11.551961
Rsp56_28 sp56_28 sp57_28 11.551961
Rsn56_28 sn56_28 sn57_28 11.551961
Rsp56_29 sp56_29 sp57_29 11.551961
Rsn56_29 sn56_29 sn57_29 11.551961
Rsp56_30 sp56_30 sp57_30 11.551961
Rsn56_30 sn56_30 sn57_30 11.551961
Rsp56_31 sp56_31 sp57_31 11.551961
Rsn56_31 sn56_31 sn57_31 11.551961
Rsp56_32 sp56_32 sp57_32 11.551961
Rsn56_32 sn56_32 sn57_32 11.551961
Rsp56_33 sp56_33 sp57_33 11.551961
Rsn56_33 sn56_33 sn57_33 11.551961
Rsp56_34 sp56_34 sp57_34 11.551961
Rsn56_34 sn56_34 sn57_34 11.551961
Rsp56_35 sp56_35 sp57_35 11.551961
Rsn56_35 sn56_35 sn57_35 11.551961
Rsp56_36 sp56_36 sp57_36 11.551961
Rsn56_36 sn56_36 sn57_36 11.551961
Rsp56_37 sp56_37 sp57_37 11.551961
Rsn56_37 sn56_37 sn57_37 11.551961
Rsp56_38 sp56_38 sp57_38 11.551961
Rsn56_38 sn56_38 sn57_38 11.551961
Rsp56_39 sp56_39 sp57_39 11.551961
Rsn56_39 sn56_39 sn57_39 11.551961
Rsp56_40 sp56_40 sp57_40 11.551961
Rsn56_40 sn56_40 sn57_40 11.551961
Rsp56_41 sp56_41 sp57_41 11.551961
Rsn56_41 sn56_41 sn57_41 11.551961
Rsp56_42 sp56_42 sp57_42 11.551961
Rsn56_42 sn56_42 sn57_42 11.551961
Rsp56_43 sp56_43 sp57_43 11.551961
Rsn56_43 sn56_43 sn57_43 11.551961
Rsp56_44 sp56_44 sp57_44 11.551961
Rsn56_44 sn56_44 sn57_44 11.551961
Rsp56_45 sp56_45 sp57_45 11.551961
Rsn56_45 sn56_45 sn57_45 11.551961
Rsp56_46 sp56_46 sp57_46 11.551961
Rsn56_46 sn56_46 sn57_46 11.551961
Rsp56_47 sp56_47 sp57_47 11.551961
Rsn56_47 sn56_47 sn57_47 11.551961
Rsp56_48 sp56_48 sp57_48 11.551961
Rsn56_48 sn56_48 sn57_48 11.551961
Rsp56_49 sp56_49 sp57_49 11.551961
Rsn56_49 sn56_49 sn57_49 11.551961
Rsp56_50 sp56_50 sp57_50 11.551961
Rsn56_50 sn56_50 sn57_50 11.551961
Rsp56_51 sp56_51 sp57_51 11.551961
Rsn56_51 sn56_51 sn57_51 11.551961
Rsp56_52 sp56_52 sp57_52 11.551961
Rsn56_52 sn56_52 sn57_52 11.551961
Rsp56_53 sp56_53 sp57_53 11.551961
Rsn56_53 sn56_53 sn57_53 11.551961
Rsp56_54 sp56_54 sp57_54 11.551961
Rsn56_54 sn56_54 sn57_54 11.551961
Rsp56_55 sp56_55 sp57_55 11.551961
Rsn56_55 sn56_55 sn57_55 11.551961
Rsp56_56 sp56_56 sp57_56 11.551961
Rsn56_56 sn56_56 sn57_56 11.551961
Rsp56_57 sp56_57 sp57_57 11.551961
Rsn56_57 sn56_57 sn57_57 11.551961
Rsp56_58 sp56_58 sp57_58 11.551961
Rsn56_58 sn56_58 sn57_58 11.551961
Rsp56_59 sp56_59 sp57_59 11.551961
Rsn56_59 sn56_59 sn57_59 11.551961
Rsp56_60 sp56_60 sp57_60 11.551961
Rsn56_60 sn56_60 sn57_60 11.551961
Rsp56_61 sp56_61 sp57_61 11.551961
Rsn56_61 sn56_61 sn57_61 11.551961
Rsp56_62 sp56_62 sp57_62 11.551961
Rsn56_62 sn56_62 sn57_62 11.551961
Rsp56_63 sp56_63 sp57_63 11.551961
Rsn56_63 sn56_63 sn57_63 11.551961
Rsp56_64 sp56_64 sp57_64 11.551961
Rsn56_64 sn56_64 sn57_64 11.551961
Rsp56_65 sp56_65 sp57_65 11.551961
Rsn56_65 sn56_65 sn57_65 11.551961
Rsp56_66 sp56_66 sp57_66 11.551961
Rsn56_66 sn56_66 sn57_66 11.551961
Rsp56_67 sp56_67 sp57_67 11.551961
Rsn56_67 sn56_67 sn57_67 11.551961
Rsp56_68 sp56_68 sp57_68 11.551961
Rsn56_68 sn56_68 sn57_68 11.551961
Rsp56_69 sp56_69 sp57_69 11.551961
Rsn56_69 sn56_69 sn57_69 11.551961
Rsp56_70 sp56_70 sp57_70 11.551961
Rsn56_70 sn56_70 sn57_70 11.551961
Rsp56_71 sp56_71 sp57_71 11.551961
Rsn56_71 sn56_71 sn57_71 11.551961
Rsp56_72 sp56_72 sp57_72 11.551961
Rsn56_72 sn56_72 sn57_72 11.551961
Rsp56_73 sp56_73 sp57_73 11.551961
Rsn56_73 sn56_73 sn57_73 11.551961
Rsp56_74 sp56_74 sp57_74 11.551961
Rsn56_74 sn56_74 sn57_74 11.551961
Rsp56_75 sp56_75 sp57_75 11.551961
Rsn56_75 sn56_75 sn57_75 11.551961
Rsp56_76 sp56_76 sp57_76 11.551961
Rsn56_76 sn56_76 sn57_76 11.551961
Rsp56_77 sp56_77 sp57_77 11.551961
Rsn56_77 sn56_77 sn57_77 11.551961
Rsp56_78 sp56_78 sp57_78 11.551961
Rsn56_78 sn56_78 sn57_78 11.551961
Rsp56_79 sp56_79 sp57_79 11.551961
Rsn56_79 sn56_79 sn57_79 11.551961
Rsp56_80 sp56_80 sp57_80 11.551961
Rsn56_80 sn56_80 sn57_80 11.551961
Rsp56_81 sp56_81 sp57_81 11.551961
Rsn56_81 sn56_81 sn57_81 11.551961
Rsp56_82 sp56_82 sp57_82 11.551961
Rsn56_82 sn56_82 sn57_82 11.551961
Rsp56_83 sp56_83 sp57_83 11.551961
Rsn56_83 sn56_83 sn57_83 11.551961
Rsp56_84 sp56_84 sp57_84 11.551961
Rsn56_84 sn56_84 sn57_84 11.551961
Rsp57_1 sp57_1 sp58_1 11.551961
Rsn57_1 sn57_1 sn58_1 11.551961
Rsp57_2 sp57_2 sp58_2 11.551961
Rsn57_2 sn57_2 sn58_2 11.551961
Rsp57_3 sp57_3 sp58_3 11.551961
Rsn57_3 sn57_3 sn58_3 11.551961
Rsp57_4 sp57_4 sp58_4 11.551961
Rsn57_4 sn57_4 sn58_4 11.551961
Rsp57_5 sp57_5 sp58_5 11.551961
Rsn57_5 sn57_5 sn58_5 11.551961
Rsp57_6 sp57_6 sp58_6 11.551961
Rsn57_6 sn57_6 sn58_6 11.551961
Rsp57_7 sp57_7 sp58_7 11.551961
Rsn57_7 sn57_7 sn58_7 11.551961
Rsp57_8 sp57_8 sp58_8 11.551961
Rsn57_8 sn57_8 sn58_8 11.551961
Rsp57_9 sp57_9 sp58_9 11.551961
Rsn57_9 sn57_9 sn58_9 11.551961
Rsp57_10 sp57_10 sp58_10 11.551961
Rsn57_10 sn57_10 sn58_10 11.551961
Rsp57_11 sp57_11 sp58_11 11.551961
Rsn57_11 sn57_11 sn58_11 11.551961
Rsp57_12 sp57_12 sp58_12 11.551961
Rsn57_12 sn57_12 sn58_12 11.551961
Rsp57_13 sp57_13 sp58_13 11.551961
Rsn57_13 sn57_13 sn58_13 11.551961
Rsp57_14 sp57_14 sp58_14 11.551961
Rsn57_14 sn57_14 sn58_14 11.551961
Rsp57_15 sp57_15 sp58_15 11.551961
Rsn57_15 sn57_15 sn58_15 11.551961
Rsp57_16 sp57_16 sp58_16 11.551961
Rsn57_16 sn57_16 sn58_16 11.551961
Rsp57_17 sp57_17 sp58_17 11.551961
Rsn57_17 sn57_17 sn58_17 11.551961
Rsp57_18 sp57_18 sp58_18 11.551961
Rsn57_18 sn57_18 sn58_18 11.551961
Rsp57_19 sp57_19 sp58_19 11.551961
Rsn57_19 sn57_19 sn58_19 11.551961
Rsp57_20 sp57_20 sp58_20 11.551961
Rsn57_20 sn57_20 sn58_20 11.551961
Rsp57_21 sp57_21 sp58_21 11.551961
Rsn57_21 sn57_21 sn58_21 11.551961
Rsp57_22 sp57_22 sp58_22 11.551961
Rsn57_22 sn57_22 sn58_22 11.551961
Rsp57_23 sp57_23 sp58_23 11.551961
Rsn57_23 sn57_23 sn58_23 11.551961
Rsp57_24 sp57_24 sp58_24 11.551961
Rsn57_24 sn57_24 sn58_24 11.551961
Rsp57_25 sp57_25 sp58_25 11.551961
Rsn57_25 sn57_25 sn58_25 11.551961
Rsp57_26 sp57_26 sp58_26 11.551961
Rsn57_26 sn57_26 sn58_26 11.551961
Rsp57_27 sp57_27 sp58_27 11.551961
Rsn57_27 sn57_27 sn58_27 11.551961
Rsp57_28 sp57_28 sp58_28 11.551961
Rsn57_28 sn57_28 sn58_28 11.551961
Rsp57_29 sp57_29 sp58_29 11.551961
Rsn57_29 sn57_29 sn58_29 11.551961
Rsp57_30 sp57_30 sp58_30 11.551961
Rsn57_30 sn57_30 sn58_30 11.551961
Rsp57_31 sp57_31 sp58_31 11.551961
Rsn57_31 sn57_31 sn58_31 11.551961
Rsp57_32 sp57_32 sp58_32 11.551961
Rsn57_32 sn57_32 sn58_32 11.551961
Rsp57_33 sp57_33 sp58_33 11.551961
Rsn57_33 sn57_33 sn58_33 11.551961
Rsp57_34 sp57_34 sp58_34 11.551961
Rsn57_34 sn57_34 sn58_34 11.551961
Rsp57_35 sp57_35 sp58_35 11.551961
Rsn57_35 sn57_35 sn58_35 11.551961
Rsp57_36 sp57_36 sp58_36 11.551961
Rsn57_36 sn57_36 sn58_36 11.551961
Rsp57_37 sp57_37 sp58_37 11.551961
Rsn57_37 sn57_37 sn58_37 11.551961
Rsp57_38 sp57_38 sp58_38 11.551961
Rsn57_38 sn57_38 sn58_38 11.551961
Rsp57_39 sp57_39 sp58_39 11.551961
Rsn57_39 sn57_39 sn58_39 11.551961
Rsp57_40 sp57_40 sp58_40 11.551961
Rsn57_40 sn57_40 sn58_40 11.551961
Rsp57_41 sp57_41 sp58_41 11.551961
Rsn57_41 sn57_41 sn58_41 11.551961
Rsp57_42 sp57_42 sp58_42 11.551961
Rsn57_42 sn57_42 sn58_42 11.551961
Rsp57_43 sp57_43 sp58_43 11.551961
Rsn57_43 sn57_43 sn58_43 11.551961
Rsp57_44 sp57_44 sp58_44 11.551961
Rsn57_44 sn57_44 sn58_44 11.551961
Rsp57_45 sp57_45 sp58_45 11.551961
Rsn57_45 sn57_45 sn58_45 11.551961
Rsp57_46 sp57_46 sp58_46 11.551961
Rsn57_46 sn57_46 sn58_46 11.551961
Rsp57_47 sp57_47 sp58_47 11.551961
Rsn57_47 sn57_47 sn58_47 11.551961
Rsp57_48 sp57_48 sp58_48 11.551961
Rsn57_48 sn57_48 sn58_48 11.551961
Rsp57_49 sp57_49 sp58_49 11.551961
Rsn57_49 sn57_49 sn58_49 11.551961
Rsp57_50 sp57_50 sp58_50 11.551961
Rsn57_50 sn57_50 sn58_50 11.551961
Rsp57_51 sp57_51 sp58_51 11.551961
Rsn57_51 sn57_51 sn58_51 11.551961
Rsp57_52 sp57_52 sp58_52 11.551961
Rsn57_52 sn57_52 sn58_52 11.551961
Rsp57_53 sp57_53 sp58_53 11.551961
Rsn57_53 sn57_53 sn58_53 11.551961
Rsp57_54 sp57_54 sp58_54 11.551961
Rsn57_54 sn57_54 sn58_54 11.551961
Rsp57_55 sp57_55 sp58_55 11.551961
Rsn57_55 sn57_55 sn58_55 11.551961
Rsp57_56 sp57_56 sp58_56 11.551961
Rsn57_56 sn57_56 sn58_56 11.551961
Rsp57_57 sp57_57 sp58_57 11.551961
Rsn57_57 sn57_57 sn58_57 11.551961
Rsp57_58 sp57_58 sp58_58 11.551961
Rsn57_58 sn57_58 sn58_58 11.551961
Rsp57_59 sp57_59 sp58_59 11.551961
Rsn57_59 sn57_59 sn58_59 11.551961
Rsp57_60 sp57_60 sp58_60 11.551961
Rsn57_60 sn57_60 sn58_60 11.551961
Rsp57_61 sp57_61 sp58_61 11.551961
Rsn57_61 sn57_61 sn58_61 11.551961
Rsp57_62 sp57_62 sp58_62 11.551961
Rsn57_62 sn57_62 sn58_62 11.551961
Rsp57_63 sp57_63 sp58_63 11.551961
Rsn57_63 sn57_63 sn58_63 11.551961
Rsp57_64 sp57_64 sp58_64 11.551961
Rsn57_64 sn57_64 sn58_64 11.551961
Rsp57_65 sp57_65 sp58_65 11.551961
Rsn57_65 sn57_65 sn58_65 11.551961
Rsp57_66 sp57_66 sp58_66 11.551961
Rsn57_66 sn57_66 sn58_66 11.551961
Rsp57_67 sp57_67 sp58_67 11.551961
Rsn57_67 sn57_67 sn58_67 11.551961
Rsp57_68 sp57_68 sp58_68 11.551961
Rsn57_68 sn57_68 sn58_68 11.551961
Rsp57_69 sp57_69 sp58_69 11.551961
Rsn57_69 sn57_69 sn58_69 11.551961
Rsp57_70 sp57_70 sp58_70 11.551961
Rsn57_70 sn57_70 sn58_70 11.551961
Rsp57_71 sp57_71 sp58_71 11.551961
Rsn57_71 sn57_71 sn58_71 11.551961
Rsp57_72 sp57_72 sp58_72 11.551961
Rsn57_72 sn57_72 sn58_72 11.551961
Rsp57_73 sp57_73 sp58_73 11.551961
Rsn57_73 sn57_73 sn58_73 11.551961
Rsp57_74 sp57_74 sp58_74 11.551961
Rsn57_74 sn57_74 sn58_74 11.551961
Rsp57_75 sp57_75 sp58_75 11.551961
Rsn57_75 sn57_75 sn58_75 11.551961
Rsp57_76 sp57_76 sp58_76 11.551961
Rsn57_76 sn57_76 sn58_76 11.551961
Rsp57_77 sp57_77 sp58_77 11.551961
Rsn57_77 sn57_77 sn58_77 11.551961
Rsp57_78 sp57_78 sp58_78 11.551961
Rsn57_78 sn57_78 sn58_78 11.551961
Rsp57_79 sp57_79 sp58_79 11.551961
Rsn57_79 sn57_79 sn58_79 11.551961
Rsp57_80 sp57_80 sp58_80 11.551961
Rsn57_80 sn57_80 sn58_80 11.551961
Rsp57_81 sp57_81 sp58_81 11.551961
Rsn57_81 sn57_81 sn58_81 11.551961
Rsp57_82 sp57_82 sp58_82 11.551961
Rsn57_82 sn57_82 sn58_82 11.551961
Rsp57_83 sp57_83 sp58_83 11.551961
Rsn57_83 sn57_83 sn58_83 11.551961
Rsp57_84 sp57_84 sp58_84 11.551961
Rsn57_84 sn57_84 sn58_84 11.551961
Rsp58_1 sp58_1 sp59_1 11.551961
Rsn58_1 sn58_1 sn59_1 11.551961
Rsp58_2 sp58_2 sp59_2 11.551961
Rsn58_2 sn58_2 sn59_2 11.551961
Rsp58_3 sp58_3 sp59_3 11.551961
Rsn58_3 sn58_3 sn59_3 11.551961
Rsp58_4 sp58_4 sp59_4 11.551961
Rsn58_4 sn58_4 sn59_4 11.551961
Rsp58_5 sp58_5 sp59_5 11.551961
Rsn58_5 sn58_5 sn59_5 11.551961
Rsp58_6 sp58_6 sp59_6 11.551961
Rsn58_6 sn58_6 sn59_6 11.551961
Rsp58_7 sp58_7 sp59_7 11.551961
Rsn58_7 sn58_7 sn59_7 11.551961
Rsp58_8 sp58_8 sp59_8 11.551961
Rsn58_8 sn58_8 sn59_8 11.551961
Rsp58_9 sp58_9 sp59_9 11.551961
Rsn58_9 sn58_9 sn59_9 11.551961
Rsp58_10 sp58_10 sp59_10 11.551961
Rsn58_10 sn58_10 sn59_10 11.551961
Rsp58_11 sp58_11 sp59_11 11.551961
Rsn58_11 sn58_11 sn59_11 11.551961
Rsp58_12 sp58_12 sp59_12 11.551961
Rsn58_12 sn58_12 sn59_12 11.551961
Rsp58_13 sp58_13 sp59_13 11.551961
Rsn58_13 sn58_13 sn59_13 11.551961
Rsp58_14 sp58_14 sp59_14 11.551961
Rsn58_14 sn58_14 sn59_14 11.551961
Rsp58_15 sp58_15 sp59_15 11.551961
Rsn58_15 sn58_15 sn59_15 11.551961
Rsp58_16 sp58_16 sp59_16 11.551961
Rsn58_16 sn58_16 sn59_16 11.551961
Rsp58_17 sp58_17 sp59_17 11.551961
Rsn58_17 sn58_17 sn59_17 11.551961
Rsp58_18 sp58_18 sp59_18 11.551961
Rsn58_18 sn58_18 sn59_18 11.551961
Rsp58_19 sp58_19 sp59_19 11.551961
Rsn58_19 sn58_19 sn59_19 11.551961
Rsp58_20 sp58_20 sp59_20 11.551961
Rsn58_20 sn58_20 sn59_20 11.551961
Rsp58_21 sp58_21 sp59_21 11.551961
Rsn58_21 sn58_21 sn59_21 11.551961
Rsp58_22 sp58_22 sp59_22 11.551961
Rsn58_22 sn58_22 sn59_22 11.551961
Rsp58_23 sp58_23 sp59_23 11.551961
Rsn58_23 sn58_23 sn59_23 11.551961
Rsp58_24 sp58_24 sp59_24 11.551961
Rsn58_24 sn58_24 sn59_24 11.551961
Rsp58_25 sp58_25 sp59_25 11.551961
Rsn58_25 sn58_25 sn59_25 11.551961
Rsp58_26 sp58_26 sp59_26 11.551961
Rsn58_26 sn58_26 sn59_26 11.551961
Rsp58_27 sp58_27 sp59_27 11.551961
Rsn58_27 sn58_27 sn59_27 11.551961
Rsp58_28 sp58_28 sp59_28 11.551961
Rsn58_28 sn58_28 sn59_28 11.551961
Rsp58_29 sp58_29 sp59_29 11.551961
Rsn58_29 sn58_29 sn59_29 11.551961
Rsp58_30 sp58_30 sp59_30 11.551961
Rsn58_30 sn58_30 sn59_30 11.551961
Rsp58_31 sp58_31 sp59_31 11.551961
Rsn58_31 sn58_31 sn59_31 11.551961
Rsp58_32 sp58_32 sp59_32 11.551961
Rsn58_32 sn58_32 sn59_32 11.551961
Rsp58_33 sp58_33 sp59_33 11.551961
Rsn58_33 sn58_33 sn59_33 11.551961
Rsp58_34 sp58_34 sp59_34 11.551961
Rsn58_34 sn58_34 sn59_34 11.551961
Rsp58_35 sp58_35 sp59_35 11.551961
Rsn58_35 sn58_35 sn59_35 11.551961
Rsp58_36 sp58_36 sp59_36 11.551961
Rsn58_36 sn58_36 sn59_36 11.551961
Rsp58_37 sp58_37 sp59_37 11.551961
Rsn58_37 sn58_37 sn59_37 11.551961
Rsp58_38 sp58_38 sp59_38 11.551961
Rsn58_38 sn58_38 sn59_38 11.551961
Rsp58_39 sp58_39 sp59_39 11.551961
Rsn58_39 sn58_39 sn59_39 11.551961
Rsp58_40 sp58_40 sp59_40 11.551961
Rsn58_40 sn58_40 sn59_40 11.551961
Rsp58_41 sp58_41 sp59_41 11.551961
Rsn58_41 sn58_41 sn59_41 11.551961
Rsp58_42 sp58_42 sp59_42 11.551961
Rsn58_42 sn58_42 sn59_42 11.551961
Rsp58_43 sp58_43 sp59_43 11.551961
Rsn58_43 sn58_43 sn59_43 11.551961
Rsp58_44 sp58_44 sp59_44 11.551961
Rsn58_44 sn58_44 sn59_44 11.551961
Rsp58_45 sp58_45 sp59_45 11.551961
Rsn58_45 sn58_45 sn59_45 11.551961
Rsp58_46 sp58_46 sp59_46 11.551961
Rsn58_46 sn58_46 sn59_46 11.551961
Rsp58_47 sp58_47 sp59_47 11.551961
Rsn58_47 sn58_47 sn59_47 11.551961
Rsp58_48 sp58_48 sp59_48 11.551961
Rsn58_48 sn58_48 sn59_48 11.551961
Rsp58_49 sp58_49 sp59_49 11.551961
Rsn58_49 sn58_49 sn59_49 11.551961
Rsp58_50 sp58_50 sp59_50 11.551961
Rsn58_50 sn58_50 sn59_50 11.551961
Rsp58_51 sp58_51 sp59_51 11.551961
Rsn58_51 sn58_51 sn59_51 11.551961
Rsp58_52 sp58_52 sp59_52 11.551961
Rsn58_52 sn58_52 sn59_52 11.551961
Rsp58_53 sp58_53 sp59_53 11.551961
Rsn58_53 sn58_53 sn59_53 11.551961
Rsp58_54 sp58_54 sp59_54 11.551961
Rsn58_54 sn58_54 sn59_54 11.551961
Rsp58_55 sp58_55 sp59_55 11.551961
Rsn58_55 sn58_55 sn59_55 11.551961
Rsp58_56 sp58_56 sp59_56 11.551961
Rsn58_56 sn58_56 sn59_56 11.551961
Rsp58_57 sp58_57 sp59_57 11.551961
Rsn58_57 sn58_57 sn59_57 11.551961
Rsp58_58 sp58_58 sp59_58 11.551961
Rsn58_58 sn58_58 sn59_58 11.551961
Rsp58_59 sp58_59 sp59_59 11.551961
Rsn58_59 sn58_59 sn59_59 11.551961
Rsp58_60 sp58_60 sp59_60 11.551961
Rsn58_60 sn58_60 sn59_60 11.551961
Rsp58_61 sp58_61 sp59_61 11.551961
Rsn58_61 sn58_61 sn59_61 11.551961
Rsp58_62 sp58_62 sp59_62 11.551961
Rsn58_62 sn58_62 sn59_62 11.551961
Rsp58_63 sp58_63 sp59_63 11.551961
Rsn58_63 sn58_63 sn59_63 11.551961
Rsp58_64 sp58_64 sp59_64 11.551961
Rsn58_64 sn58_64 sn59_64 11.551961
Rsp58_65 sp58_65 sp59_65 11.551961
Rsn58_65 sn58_65 sn59_65 11.551961
Rsp58_66 sp58_66 sp59_66 11.551961
Rsn58_66 sn58_66 sn59_66 11.551961
Rsp58_67 sp58_67 sp59_67 11.551961
Rsn58_67 sn58_67 sn59_67 11.551961
Rsp58_68 sp58_68 sp59_68 11.551961
Rsn58_68 sn58_68 sn59_68 11.551961
Rsp58_69 sp58_69 sp59_69 11.551961
Rsn58_69 sn58_69 sn59_69 11.551961
Rsp58_70 sp58_70 sp59_70 11.551961
Rsn58_70 sn58_70 sn59_70 11.551961
Rsp58_71 sp58_71 sp59_71 11.551961
Rsn58_71 sn58_71 sn59_71 11.551961
Rsp58_72 sp58_72 sp59_72 11.551961
Rsn58_72 sn58_72 sn59_72 11.551961
Rsp58_73 sp58_73 sp59_73 11.551961
Rsn58_73 sn58_73 sn59_73 11.551961
Rsp58_74 sp58_74 sp59_74 11.551961
Rsn58_74 sn58_74 sn59_74 11.551961
Rsp58_75 sp58_75 sp59_75 11.551961
Rsn58_75 sn58_75 sn59_75 11.551961
Rsp58_76 sp58_76 sp59_76 11.551961
Rsn58_76 sn58_76 sn59_76 11.551961
Rsp58_77 sp58_77 sp59_77 11.551961
Rsn58_77 sn58_77 sn59_77 11.551961
Rsp58_78 sp58_78 sp59_78 11.551961
Rsn58_78 sn58_78 sn59_78 11.551961
Rsp58_79 sp58_79 sp59_79 11.551961
Rsn58_79 sn58_79 sn59_79 11.551961
Rsp58_80 sp58_80 sp59_80 11.551961
Rsn58_80 sn58_80 sn59_80 11.551961
Rsp58_81 sp58_81 sp59_81 11.551961
Rsn58_81 sn58_81 sn59_81 11.551961
Rsp58_82 sp58_82 sp59_82 11.551961
Rsn58_82 sn58_82 sn59_82 11.551961
Rsp58_83 sp58_83 sp59_83 11.551961
Rsn58_83 sn58_83 sn59_83 11.551961
Rsp58_84 sp58_84 sp59_84 11.551961
Rsn58_84 sn58_84 sn59_84 11.551961
Rsp59_1 sp59_1 sp60_1 11.551961
Rsn59_1 sn59_1 sn60_1 11.551961
Rsp59_2 sp59_2 sp60_2 11.551961
Rsn59_2 sn59_2 sn60_2 11.551961
Rsp59_3 sp59_3 sp60_3 11.551961
Rsn59_3 sn59_3 sn60_3 11.551961
Rsp59_4 sp59_4 sp60_4 11.551961
Rsn59_4 sn59_4 sn60_4 11.551961
Rsp59_5 sp59_5 sp60_5 11.551961
Rsn59_5 sn59_5 sn60_5 11.551961
Rsp59_6 sp59_6 sp60_6 11.551961
Rsn59_6 sn59_6 sn60_6 11.551961
Rsp59_7 sp59_7 sp60_7 11.551961
Rsn59_7 sn59_7 sn60_7 11.551961
Rsp59_8 sp59_8 sp60_8 11.551961
Rsn59_8 sn59_8 sn60_8 11.551961
Rsp59_9 sp59_9 sp60_9 11.551961
Rsn59_9 sn59_9 sn60_9 11.551961
Rsp59_10 sp59_10 sp60_10 11.551961
Rsn59_10 sn59_10 sn60_10 11.551961
Rsp59_11 sp59_11 sp60_11 11.551961
Rsn59_11 sn59_11 sn60_11 11.551961
Rsp59_12 sp59_12 sp60_12 11.551961
Rsn59_12 sn59_12 sn60_12 11.551961
Rsp59_13 sp59_13 sp60_13 11.551961
Rsn59_13 sn59_13 sn60_13 11.551961
Rsp59_14 sp59_14 sp60_14 11.551961
Rsn59_14 sn59_14 sn60_14 11.551961
Rsp59_15 sp59_15 sp60_15 11.551961
Rsn59_15 sn59_15 sn60_15 11.551961
Rsp59_16 sp59_16 sp60_16 11.551961
Rsn59_16 sn59_16 sn60_16 11.551961
Rsp59_17 sp59_17 sp60_17 11.551961
Rsn59_17 sn59_17 sn60_17 11.551961
Rsp59_18 sp59_18 sp60_18 11.551961
Rsn59_18 sn59_18 sn60_18 11.551961
Rsp59_19 sp59_19 sp60_19 11.551961
Rsn59_19 sn59_19 sn60_19 11.551961
Rsp59_20 sp59_20 sp60_20 11.551961
Rsn59_20 sn59_20 sn60_20 11.551961
Rsp59_21 sp59_21 sp60_21 11.551961
Rsn59_21 sn59_21 sn60_21 11.551961
Rsp59_22 sp59_22 sp60_22 11.551961
Rsn59_22 sn59_22 sn60_22 11.551961
Rsp59_23 sp59_23 sp60_23 11.551961
Rsn59_23 sn59_23 sn60_23 11.551961
Rsp59_24 sp59_24 sp60_24 11.551961
Rsn59_24 sn59_24 sn60_24 11.551961
Rsp59_25 sp59_25 sp60_25 11.551961
Rsn59_25 sn59_25 sn60_25 11.551961
Rsp59_26 sp59_26 sp60_26 11.551961
Rsn59_26 sn59_26 sn60_26 11.551961
Rsp59_27 sp59_27 sp60_27 11.551961
Rsn59_27 sn59_27 sn60_27 11.551961
Rsp59_28 sp59_28 sp60_28 11.551961
Rsn59_28 sn59_28 sn60_28 11.551961
Rsp59_29 sp59_29 sp60_29 11.551961
Rsn59_29 sn59_29 sn60_29 11.551961
Rsp59_30 sp59_30 sp60_30 11.551961
Rsn59_30 sn59_30 sn60_30 11.551961
Rsp59_31 sp59_31 sp60_31 11.551961
Rsn59_31 sn59_31 sn60_31 11.551961
Rsp59_32 sp59_32 sp60_32 11.551961
Rsn59_32 sn59_32 sn60_32 11.551961
Rsp59_33 sp59_33 sp60_33 11.551961
Rsn59_33 sn59_33 sn60_33 11.551961
Rsp59_34 sp59_34 sp60_34 11.551961
Rsn59_34 sn59_34 sn60_34 11.551961
Rsp59_35 sp59_35 sp60_35 11.551961
Rsn59_35 sn59_35 sn60_35 11.551961
Rsp59_36 sp59_36 sp60_36 11.551961
Rsn59_36 sn59_36 sn60_36 11.551961
Rsp59_37 sp59_37 sp60_37 11.551961
Rsn59_37 sn59_37 sn60_37 11.551961
Rsp59_38 sp59_38 sp60_38 11.551961
Rsn59_38 sn59_38 sn60_38 11.551961
Rsp59_39 sp59_39 sp60_39 11.551961
Rsn59_39 sn59_39 sn60_39 11.551961
Rsp59_40 sp59_40 sp60_40 11.551961
Rsn59_40 sn59_40 sn60_40 11.551961
Rsp59_41 sp59_41 sp60_41 11.551961
Rsn59_41 sn59_41 sn60_41 11.551961
Rsp59_42 sp59_42 sp60_42 11.551961
Rsn59_42 sn59_42 sn60_42 11.551961
Rsp59_43 sp59_43 sp60_43 11.551961
Rsn59_43 sn59_43 sn60_43 11.551961
Rsp59_44 sp59_44 sp60_44 11.551961
Rsn59_44 sn59_44 sn60_44 11.551961
Rsp59_45 sp59_45 sp60_45 11.551961
Rsn59_45 sn59_45 sn60_45 11.551961
Rsp59_46 sp59_46 sp60_46 11.551961
Rsn59_46 sn59_46 sn60_46 11.551961
Rsp59_47 sp59_47 sp60_47 11.551961
Rsn59_47 sn59_47 sn60_47 11.551961
Rsp59_48 sp59_48 sp60_48 11.551961
Rsn59_48 sn59_48 sn60_48 11.551961
Rsp59_49 sp59_49 sp60_49 11.551961
Rsn59_49 sn59_49 sn60_49 11.551961
Rsp59_50 sp59_50 sp60_50 11.551961
Rsn59_50 sn59_50 sn60_50 11.551961
Rsp59_51 sp59_51 sp60_51 11.551961
Rsn59_51 sn59_51 sn60_51 11.551961
Rsp59_52 sp59_52 sp60_52 11.551961
Rsn59_52 sn59_52 sn60_52 11.551961
Rsp59_53 sp59_53 sp60_53 11.551961
Rsn59_53 sn59_53 sn60_53 11.551961
Rsp59_54 sp59_54 sp60_54 11.551961
Rsn59_54 sn59_54 sn60_54 11.551961
Rsp59_55 sp59_55 sp60_55 11.551961
Rsn59_55 sn59_55 sn60_55 11.551961
Rsp59_56 sp59_56 sp60_56 11.551961
Rsn59_56 sn59_56 sn60_56 11.551961
Rsp59_57 sp59_57 sp60_57 11.551961
Rsn59_57 sn59_57 sn60_57 11.551961
Rsp59_58 sp59_58 sp60_58 11.551961
Rsn59_58 sn59_58 sn60_58 11.551961
Rsp59_59 sp59_59 sp60_59 11.551961
Rsn59_59 sn59_59 sn60_59 11.551961
Rsp59_60 sp59_60 sp60_60 11.551961
Rsn59_60 sn59_60 sn60_60 11.551961
Rsp59_61 sp59_61 sp60_61 11.551961
Rsn59_61 sn59_61 sn60_61 11.551961
Rsp59_62 sp59_62 sp60_62 11.551961
Rsn59_62 sn59_62 sn60_62 11.551961
Rsp59_63 sp59_63 sp60_63 11.551961
Rsn59_63 sn59_63 sn60_63 11.551961
Rsp59_64 sp59_64 sp60_64 11.551961
Rsn59_64 sn59_64 sn60_64 11.551961
Rsp59_65 sp59_65 sp60_65 11.551961
Rsn59_65 sn59_65 sn60_65 11.551961
Rsp59_66 sp59_66 sp60_66 11.551961
Rsn59_66 sn59_66 sn60_66 11.551961
Rsp59_67 sp59_67 sp60_67 11.551961
Rsn59_67 sn59_67 sn60_67 11.551961
Rsp59_68 sp59_68 sp60_68 11.551961
Rsn59_68 sn59_68 sn60_68 11.551961
Rsp59_69 sp59_69 sp60_69 11.551961
Rsn59_69 sn59_69 sn60_69 11.551961
Rsp59_70 sp59_70 sp60_70 11.551961
Rsn59_70 sn59_70 sn60_70 11.551961
Rsp59_71 sp59_71 sp60_71 11.551961
Rsn59_71 sn59_71 sn60_71 11.551961
Rsp59_72 sp59_72 sp60_72 11.551961
Rsn59_72 sn59_72 sn60_72 11.551961
Rsp59_73 sp59_73 sp60_73 11.551961
Rsn59_73 sn59_73 sn60_73 11.551961
Rsp59_74 sp59_74 sp60_74 11.551961
Rsn59_74 sn59_74 sn60_74 11.551961
Rsp59_75 sp59_75 sp60_75 11.551961
Rsn59_75 sn59_75 sn60_75 11.551961
Rsp59_76 sp59_76 sp60_76 11.551961
Rsn59_76 sn59_76 sn60_76 11.551961
Rsp59_77 sp59_77 sp60_77 11.551961
Rsn59_77 sn59_77 sn60_77 11.551961
Rsp59_78 sp59_78 sp60_78 11.551961
Rsn59_78 sn59_78 sn60_78 11.551961
Rsp59_79 sp59_79 sp60_79 11.551961
Rsn59_79 sn59_79 sn60_79 11.551961
Rsp59_80 sp59_80 sp60_80 11.551961
Rsn59_80 sn59_80 sn60_80 11.551961
Rsp59_81 sp59_81 sp60_81 11.551961
Rsn59_81 sn59_81 sn60_81 11.551961
Rsp59_82 sp59_82 sp60_82 11.551961
Rsn59_82 sn59_82 sn60_82 11.551961
Rsp59_83 sp59_83 sp60_83 11.551961
Rsn59_83 sn59_83 sn60_83 11.551961
Rsp59_84 sp59_84 sp60_84 11.551961
Rsn59_84 sn59_84 sn60_84 11.551961
Rsp60_1 sp60_1 sp61_1 11.551961
Rsn60_1 sn60_1 sn61_1 11.551961
Rsp60_2 sp60_2 sp61_2 11.551961
Rsn60_2 sn60_2 sn61_2 11.551961
Rsp60_3 sp60_3 sp61_3 11.551961
Rsn60_3 sn60_3 sn61_3 11.551961
Rsp60_4 sp60_4 sp61_4 11.551961
Rsn60_4 sn60_4 sn61_4 11.551961
Rsp60_5 sp60_5 sp61_5 11.551961
Rsn60_5 sn60_5 sn61_5 11.551961
Rsp60_6 sp60_6 sp61_6 11.551961
Rsn60_6 sn60_6 sn61_6 11.551961
Rsp60_7 sp60_7 sp61_7 11.551961
Rsn60_7 sn60_7 sn61_7 11.551961
Rsp60_8 sp60_8 sp61_8 11.551961
Rsn60_8 sn60_8 sn61_8 11.551961
Rsp60_9 sp60_9 sp61_9 11.551961
Rsn60_9 sn60_9 sn61_9 11.551961
Rsp60_10 sp60_10 sp61_10 11.551961
Rsn60_10 sn60_10 sn61_10 11.551961
Rsp60_11 sp60_11 sp61_11 11.551961
Rsn60_11 sn60_11 sn61_11 11.551961
Rsp60_12 sp60_12 sp61_12 11.551961
Rsn60_12 sn60_12 sn61_12 11.551961
Rsp60_13 sp60_13 sp61_13 11.551961
Rsn60_13 sn60_13 sn61_13 11.551961
Rsp60_14 sp60_14 sp61_14 11.551961
Rsn60_14 sn60_14 sn61_14 11.551961
Rsp60_15 sp60_15 sp61_15 11.551961
Rsn60_15 sn60_15 sn61_15 11.551961
Rsp60_16 sp60_16 sp61_16 11.551961
Rsn60_16 sn60_16 sn61_16 11.551961
Rsp60_17 sp60_17 sp61_17 11.551961
Rsn60_17 sn60_17 sn61_17 11.551961
Rsp60_18 sp60_18 sp61_18 11.551961
Rsn60_18 sn60_18 sn61_18 11.551961
Rsp60_19 sp60_19 sp61_19 11.551961
Rsn60_19 sn60_19 sn61_19 11.551961
Rsp60_20 sp60_20 sp61_20 11.551961
Rsn60_20 sn60_20 sn61_20 11.551961
Rsp60_21 sp60_21 sp61_21 11.551961
Rsn60_21 sn60_21 sn61_21 11.551961
Rsp60_22 sp60_22 sp61_22 11.551961
Rsn60_22 sn60_22 sn61_22 11.551961
Rsp60_23 sp60_23 sp61_23 11.551961
Rsn60_23 sn60_23 sn61_23 11.551961
Rsp60_24 sp60_24 sp61_24 11.551961
Rsn60_24 sn60_24 sn61_24 11.551961
Rsp60_25 sp60_25 sp61_25 11.551961
Rsn60_25 sn60_25 sn61_25 11.551961
Rsp60_26 sp60_26 sp61_26 11.551961
Rsn60_26 sn60_26 sn61_26 11.551961
Rsp60_27 sp60_27 sp61_27 11.551961
Rsn60_27 sn60_27 sn61_27 11.551961
Rsp60_28 sp60_28 sp61_28 11.551961
Rsn60_28 sn60_28 sn61_28 11.551961
Rsp60_29 sp60_29 sp61_29 11.551961
Rsn60_29 sn60_29 sn61_29 11.551961
Rsp60_30 sp60_30 sp61_30 11.551961
Rsn60_30 sn60_30 sn61_30 11.551961
Rsp60_31 sp60_31 sp61_31 11.551961
Rsn60_31 sn60_31 sn61_31 11.551961
Rsp60_32 sp60_32 sp61_32 11.551961
Rsn60_32 sn60_32 sn61_32 11.551961
Rsp60_33 sp60_33 sp61_33 11.551961
Rsn60_33 sn60_33 sn61_33 11.551961
Rsp60_34 sp60_34 sp61_34 11.551961
Rsn60_34 sn60_34 sn61_34 11.551961
Rsp60_35 sp60_35 sp61_35 11.551961
Rsn60_35 sn60_35 sn61_35 11.551961
Rsp60_36 sp60_36 sp61_36 11.551961
Rsn60_36 sn60_36 sn61_36 11.551961
Rsp60_37 sp60_37 sp61_37 11.551961
Rsn60_37 sn60_37 sn61_37 11.551961
Rsp60_38 sp60_38 sp61_38 11.551961
Rsn60_38 sn60_38 sn61_38 11.551961
Rsp60_39 sp60_39 sp61_39 11.551961
Rsn60_39 sn60_39 sn61_39 11.551961
Rsp60_40 sp60_40 sp61_40 11.551961
Rsn60_40 sn60_40 sn61_40 11.551961
Rsp60_41 sp60_41 sp61_41 11.551961
Rsn60_41 sn60_41 sn61_41 11.551961
Rsp60_42 sp60_42 sp61_42 11.551961
Rsn60_42 sn60_42 sn61_42 11.551961
Rsp60_43 sp60_43 sp61_43 11.551961
Rsn60_43 sn60_43 sn61_43 11.551961
Rsp60_44 sp60_44 sp61_44 11.551961
Rsn60_44 sn60_44 sn61_44 11.551961
Rsp60_45 sp60_45 sp61_45 11.551961
Rsn60_45 sn60_45 sn61_45 11.551961
Rsp60_46 sp60_46 sp61_46 11.551961
Rsn60_46 sn60_46 sn61_46 11.551961
Rsp60_47 sp60_47 sp61_47 11.551961
Rsn60_47 sn60_47 sn61_47 11.551961
Rsp60_48 sp60_48 sp61_48 11.551961
Rsn60_48 sn60_48 sn61_48 11.551961
Rsp60_49 sp60_49 sp61_49 11.551961
Rsn60_49 sn60_49 sn61_49 11.551961
Rsp60_50 sp60_50 sp61_50 11.551961
Rsn60_50 sn60_50 sn61_50 11.551961
Rsp60_51 sp60_51 sp61_51 11.551961
Rsn60_51 sn60_51 sn61_51 11.551961
Rsp60_52 sp60_52 sp61_52 11.551961
Rsn60_52 sn60_52 sn61_52 11.551961
Rsp60_53 sp60_53 sp61_53 11.551961
Rsn60_53 sn60_53 sn61_53 11.551961
Rsp60_54 sp60_54 sp61_54 11.551961
Rsn60_54 sn60_54 sn61_54 11.551961
Rsp60_55 sp60_55 sp61_55 11.551961
Rsn60_55 sn60_55 sn61_55 11.551961
Rsp60_56 sp60_56 sp61_56 11.551961
Rsn60_56 sn60_56 sn61_56 11.551961
Rsp60_57 sp60_57 sp61_57 11.551961
Rsn60_57 sn60_57 sn61_57 11.551961
Rsp60_58 sp60_58 sp61_58 11.551961
Rsn60_58 sn60_58 sn61_58 11.551961
Rsp60_59 sp60_59 sp61_59 11.551961
Rsn60_59 sn60_59 sn61_59 11.551961
Rsp60_60 sp60_60 sp61_60 11.551961
Rsn60_60 sn60_60 sn61_60 11.551961
Rsp60_61 sp60_61 sp61_61 11.551961
Rsn60_61 sn60_61 sn61_61 11.551961
Rsp60_62 sp60_62 sp61_62 11.551961
Rsn60_62 sn60_62 sn61_62 11.551961
Rsp60_63 sp60_63 sp61_63 11.551961
Rsn60_63 sn60_63 sn61_63 11.551961
Rsp60_64 sp60_64 sp61_64 11.551961
Rsn60_64 sn60_64 sn61_64 11.551961
Rsp60_65 sp60_65 sp61_65 11.551961
Rsn60_65 sn60_65 sn61_65 11.551961
Rsp60_66 sp60_66 sp61_66 11.551961
Rsn60_66 sn60_66 sn61_66 11.551961
Rsp60_67 sp60_67 sp61_67 11.551961
Rsn60_67 sn60_67 sn61_67 11.551961
Rsp60_68 sp60_68 sp61_68 11.551961
Rsn60_68 sn60_68 sn61_68 11.551961
Rsp60_69 sp60_69 sp61_69 11.551961
Rsn60_69 sn60_69 sn61_69 11.551961
Rsp60_70 sp60_70 sp61_70 11.551961
Rsn60_70 sn60_70 sn61_70 11.551961
Rsp60_71 sp60_71 sp61_71 11.551961
Rsn60_71 sn60_71 sn61_71 11.551961
Rsp60_72 sp60_72 sp61_72 11.551961
Rsn60_72 sn60_72 sn61_72 11.551961
Rsp60_73 sp60_73 sp61_73 11.551961
Rsn60_73 sn60_73 sn61_73 11.551961
Rsp60_74 sp60_74 sp61_74 11.551961
Rsn60_74 sn60_74 sn61_74 11.551961
Rsp60_75 sp60_75 sp61_75 11.551961
Rsn60_75 sn60_75 sn61_75 11.551961
Rsp60_76 sp60_76 sp61_76 11.551961
Rsn60_76 sn60_76 sn61_76 11.551961
Rsp60_77 sp60_77 sp61_77 11.551961
Rsn60_77 sn60_77 sn61_77 11.551961
Rsp60_78 sp60_78 sp61_78 11.551961
Rsn60_78 sn60_78 sn61_78 11.551961
Rsp60_79 sp60_79 sp61_79 11.551961
Rsn60_79 sn60_79 sn61_79 11.551961
Rsp60_80 sp60_80 sp61_80 11.551961
Rsn60_80 sn60_80 sn61_80 11.551961
Rsp60_81 sp60_81 sp61_81 11.551961
Rsn60_81 sn60_81 sn61_81 11.551961
Rsp60_82 sp60_82 sp61_82 11.551961
Rsn60_82 sn60_82 sn61_82 11.551961
Rsp60_83 sp60_83 sp61_83 11.551961
Rsn60_83 sn60_83 sn61_83 11.551961
Rsp60_84 sp60_84 sp61_84 11.551961
Rsn60_84 sn60_84 sn61_84 11.551961
Rsp61_1 sp61_1 sp1_p2 11.551961
Rsn61_1 sn61_1 sn1_p2 11.551961
Rsp61_2 sp61_2 sp2_p2 11.551961
Rsn61_2 sn61_2 sn2_p2 11.551961
Rsp61_3 sp61_3 sp3_p2 11.551961
Rsn61_3 sn61_3 sn3_p2 11.551961
Rsp61_4 sp61_4 sp4_p2 11.551961
Rsn61_4 sn61_4 sn4_p2 11.551961
Rsp61_5 sp61_5 sp5_p2 11.551961
Rsn61_5 sn61_5 sn5_p2 11.551961
Rsp61_6 sp61_6 sp6_p2 11.551961
Rsn61_6 sn61_6 sn6_p2 11.551961
Rsp61_7 sp61_7 sp7_p2 11.551961
Rsn61_7 sn61_7 sn7_p2 11.551961
Rsp61_8 sp61_8 sp8_p2 11.551961
Rsn61_8 sn61_8 sn8_p2 11.551961
Rsp61_9 sp61_9 sp9_p2 11.551961
Rsn61_9 sn61_9 sn9_p2 11.551961
Rsp61_10 sp61_10 sp10_p2 11.551961
Rsn61_10 sn61_10 sn10_p2 11.551961
Rsp61_11 sp61_11 sp11_p2 11.551961
Rsn61_11 sn61_11 sn11_p2 11.551961
Rsp61_12 sp61_12 sp12_p2 11.551961
Rsn61_12 sn61_12 sn12_p2 11.551961
Rsp61_13 sp61_13 sp13_p2 11.551961
Rsn61_13 sn61_13 sn13_p2 11.551961
Rsp61_14 sp61_14 sp14_p2 11.551961
Rsn61_14 sn61_14 sn14_p2 11.551961
Rsp61_15 sp61_15 sp15_p2 11.551961
Rsn61_15 sn61_15 sn15_p2 11.551961
Rsp61_16 sp61_16 sp16_p2 11.551961
Rsn61_16 sn61_16 sn16_p2 11.551961
Rsp61_17 sp61_17 sp17_p2 11.551961
Rsn61_17 sn61_17 sn17_p2 11.551961
Rsp61_18 sp61_18 sp18_p2 11.551961
Rsn61_18 sn61_18 sn18_p2 11.551961
Rsp61_19 sp61_19 sp19_p2 11.551961
Rsn61_19 sn61_19 sn19_p2 11.551961
Rsp61_20 sp61_20 sp20_p2 11.551961
Rsn61_20 sn61_20 sn20_p2 11.551961
Rsp61_21 sp61_21 sp21_p2 11.551961
Rsn61_21 sn61_21 sn21_p2 11.551961
Rsp61_22 sp61_22 sp22_p2 11.551961
Rsn61_22 sn61_22 sn22_p2 11.551961
Rsp61_23 sp61_23 sp23_p2 11.551961
Rsn61_23 sn61_23 sn23_p2 11.551961
Rsp61_24 sp61_24 sp24_p2 11.551961
Rsn61_24 sn61_24 sn24_p2 11.551961
Rsp61_25 sp61_25 sp25_p2 11.551961
Rsn61_25 sn61_25 sn25_p2 11.551961
Rsp61_26 sp61_26 sp26_p2 11.551961
Rsn61_26 sn61_26 sn26_p2 11.551961
Rsp61_27 sp61_27 sp27_p2 11.551961
Rsn61_27 sn61_27 sn27_p2 11.551961
Rsp61_28 sp61_28 sp28_p2 11.551961
Rsn61_28 sn61_28 sn28_p2 11.551961
Rsp61_29 sp61_29 sp29_p2 11.551961
Rsn61_29 sn61_29 sn29_p2 11.551961
Rsp61_30 sp61_30 sp30_p2 11.551961
Rsn61_30 sn61_30 sn30_p2 11.551961
Rsp61_31 sp61_31 sp31_p2 11.551961
Rsn61_31 sn61_31 sn31_p2 11.551961
Rsp61_32 sp61_32 sp32_p2 11.551961
Rsn61_32 sn61_32 sn32_p2 11.551961
Rsp61_33 sp61_33 sp33_p2 11.551961
Rsn61_33 sn61_33 sn33_p2 11.551961
Rsp61_34 sp61_34 sp34_p2 11.551961
Rsn61_34 sn61_34 sn34_p2 11.551961
Rsp61_35 sp61_35 sp35_p2 11.551961
Rsn61_35 sn61_35 sn35_p2 11.551961
Rsp61_36 sp61_36 sp36_p2 11.551961
Rsn61_36 sn61_36 sn36_p2 11.551961
Rsp61_37 sp61_37 sp37_p2 11.551961
Rsn61_37 sn61_37 sn37_p2 11.551961
Rsp61_38 sp61_38 sp38_p2 11.551961
Rsn61_38 sn61_38 sn38_p2 11.551961
Rsp61_39 sp61_39 sp39_p2 11.551961
Rsn61_39 sn61_39 sn39_p2 11.551961
Rsp61_40 sp61_40 sp40_p2 11.551961
Rsn61_40 sn61_40 sn40_p2 11.551961
Rsp61_41 sp61_41 sp41_p2 11.551961
Rsn61_41 sn61_41 sn41_p2 11.551961
Rsp61_42 sp61_42 sp42_p2 11.551961
Rsn61_42 sn61_42 sn42_p2 11.551961
Rsp61_43 sp61_43 sp43_p2 11.551961
Rsn61_43 sn61_43 sn43_p2 11.551961
Rsp61_44 sp61_44 sp44_p2 11.551961
Rsn61_44 sn61_44 sn44_p2 11.551961
Rsp61_45 sp61_45 sp45_p2 11.551961
Rsn61_45 sn61_45 sn45_p2 11.551961
Rsp61_46 sp61_46 sp46_p2 11.551961
Rsn61_46 sn61_46 sn46_p2 11.551961
Rsp61_47 sp61_47 sp47_p2 11.551961
Rsn61_47 sn61_47 sn47_p2 11.551961
Rsp61_48 sp61_48 sp48_p2 11.551961
Rsn61_48 sn61_48 sn48_p2 11.551961
Rsp61_49 sp61_49 sp49_p2 11.551961
Rsn61_49 sn61_49 sn49_p2 11.551961
Rsp61_50 sp61_50 sp50_p2 11.551961
Rsn61_50 sn61_50 sn50_p2 11.551961
Rsp61_51 sp61_51 sp51_p2 11.551961
Rsn61_51 sn61_51 sn51_p2 11.551961
Rsp61_52 sp61_52 sp52_p2 11.551961
Rsn61_52 sn61_52 sn52_p2 11.551961
Rsp61_53 sp61_53 sp53_p2 11.551961
Rsn61_53 sn61_53 sn53_p2 11.551961
Rsp61_54 sp61_54 sp54_p2 11.551961
Rsn61_54 sn61_54 sn54_p2 11.551961
Rsp61_55 sp61_55 sp55_p2 11.551961
Rsn61_55 sn61_55 sn55_p2 11.551961
Rsp61_56 sp61_56 sp56_p2 11.551961
Rsn61_56 sn61_56 sn56_p2 11.551961
Rsp61_57 sp61_57 sp57_p2 11.551961
Rsn61_57 sn61_57 sn57_p2 11.551961
Rsp61_58 sp61_58 sp58_p2 11.551961
Rsn61_58 sn61_58 sn58_p2 11.551961
Rsp61_59 sp61_59 sp59_p2 11.551961
Rsn61_59 sn61_59 sn59_p2 11.551961
Rsp61_60 sp61_60 sp60_p2 11.551961
Rsn61_60 sn61_60 sn60_p2 11.551961
Rsp61_61 sp61_61 sp61_p2 11.551961
Rsn61_61 sn61_61 sn61_p2 11.551961
Rsp61_62 sp61_62 sp62_p2 11.551961
Rsn61_62 sn61_62 sn62_p2 11.551961
Rsp61_63 sp61_63 sp63_p2 11.551961
Rsn61_63 sn61_63 sn63_p2 11.551961
Rsp61_64 sp61_64 sp64_p2 11.551961
Rsn61_64 sn61_64 sn64_p2 11.551961
Rsp61_65 sp61_65 sp65_p2 11.551961
Rsn61_65 sn61_65 sn65_p2 11.551961
Rsp61_66 sp61_66 sp66_p2 11.551961
Rsn61_66 sn61_66 sn66_p2 11.551961
Rsp61_67 sp61_67 sp67_p2 11.551961
Rsn61_67 sn61_67 sn67_p2 11.551961
Rsp61_68 sp61_68 sp68_p2 11.551961
Rsn61_68 sn61_68 sn68_p2 11.551961
Rsp61_69 sp61_69 sp69_p2 11.551961
Rsn61_69 sn61_69 sn69_p2 11.551961
Rsp61_70 sp61_70 sp70_p2 11.551961
Rsn61_70 sn61_70 sn70_p2 11.551961
Rsp61_71 sp61_71 sp71_p2 11.551961
Rsn61_71 sn61_71 sn71_p2 11.551961
Rsp61_72 sp61_72 sp72_p2 11.551961
Rsn61_72 sn61_72 sn72_p2 11.551961
Rsp61_73 sp61_73 sp73_p2 11.551961
Rsn61_73 sn61_73 sn73_p2 11.551961
Rsp61_74 sp61_74 sp74_p2 11.551961
Rsn61_74 sn61_74 sn74_p2 11.551961
Rsp61_75 sp61_75 sp75_p2 11.551961
Rsn61_75 sn61_75 sn75_p2 11.551961
Rsp61_76 sp61_76 sp76_p2 11.551961
Rsn61_76 sn61_76 sn76_p2 11.551961
Rsp61_77 sp61_77 sp77_p2 11.551961
Rsn61_77 sn61_77 sn77_p2 11.551961
Rsp61_78 sp61_78 sp78_p2 11.551961
Rsn61_78 sn61_78 sn78_p2 11.551961
Rsp61_79 sp61_79 sp79_p2 11.551961
Rsn61_79 sn61_79 sn79_p2 11.551961
Rsp61_80 sp61_80 sp80_p2 11.551961
Rsn61_80 sn61_80 sn80_p2 11.551961
Rsp61_81 sp61_81 sp81_p2 11.551961
Rsn61_81 sn61_81 sn81_p2 11.551961
Rsp61_82 sp61_82 sp82_p2 11.551961
Rsn61_82 sn61_82 sn82_p2 11.551961
Rsp61_83 sp61_83 sp83_p2 11.551961
Rsn61_83 sn61_83 sn83_p2 11.551961
Rsp61_84 sp61_84 sp84_p2 11.551961
Rsn61_84 sn61_84 sn84_p2 11.551961
Rsp62_1 sp62_1 sp63_1 11.551961
Rsn62_1 sn62_1 sn63_1 11.551961
Rsp62_2 sp62_2 sp63_2 11.551961
Rsn62_2 sn62_2 sn63_2 11.551961
Rsp62_3 sp62_3 sp63_3 11.551961
Rsn62_3 sn62_3 sn63_3 11.551961
Rsp62_4 sp62_4 sp63_4 11.551961
Rsn62_4 sn62_4 sn63_4 11.551961
Rsp62_5 sp62_5 sp63_5 11.551961
Rsn62_5 sn62_5 sn63_5 11.551961
Rsp62_6 sp62_6 sp63_6 11.551961
Rsn62_6 sn62_6 sn63_6 11.551961
Rsp62_7 sp62_7 sp63_7 11.551961
Rsn62_7 sn62_7 sn63_7 11.551961
Rsp62_8 sp62_8 sp63_8 11.551961
Rsn62_8 sn62_8 sn63_8 11.551961
Rsp62_9 sp62_9 sp63_9 11.551961
Rsn62_9 sn62_9 sn63_9 11.551961
Rsp62_10 sp62_10 sp63_10 11.551961
Rsn62_10 sn62_10 sn63_10 11.551961
Rsp62_11 sp62_11 sp63_11 11.551961
Rsn62_11 sn62_11 sn63_11 11.551961
Rsp62_12 sp62_12 sp63_12 11.551961
Rsn62_12 sn62_12 sn63_12 11.551961
Rsp62_13 sp62_13 sp63_13 11.551961
Rsn62_13 sn62_13 sn63_13 11.551961
Rsp62_14 sp62_14 sp63_14 11.551961
Rsn62_14 sn62_14 sn63_14 11.551961
Rsp62_15 sp62_15 sp63_15 11.551961
Rsn62_15 sn62_15 sn63_15 11.551961
Rsp62_16 sp62_16 sp63_16 11.551961
Rsn62_16 sn62_16 sn63_16 11.551961
Rsp62_17 sp62_17 sp63_17 11.551961
Rsn62_17 sn62_17 sn63_17 11.551961
Rsp62_18 sp62_18 sp63_18 11.551961
Rsn62_18 sn62_18 sn63_18 11.551961
Rsp62_19 sp62_19 sp63_19 11.551961
Rsn62_19 sn62_19 sn63_19 11.551961
Rsp62_20 sp62_20 sp63_20 11.551961
Rsn62_20 sn62_20 sn63_20 11.551961
Rsp62_21 sp62_21 sp63_21 11.551961
Rsn62_21 sn62_21 sn63_21 11.551961
Rsp62_22 sp62_22 sp63_22 11.551961
Rsn62_22 sn62_22 sn63_22 11.551961
Rsp62_23 sp62_23 sp63_23 11.551961
Rsn62_23 sn62_23 sn63_23 11.551961
Rsp62_24 sp62_24 sp63_24 11.551961
Rsn62_24 sn62_24 sn63_24 11.551961
Rsp62_25 sp62_25 sp63_25 11.551961
Rsn62_25 sn62_25 sn63_25 11.551961
Rsp62_26 sp62_26 sp63_26 11.551961
Rsn62_26 sn62_26 sn63_26 11.551961
Rsp62_27 sp62_27 sp63_27 11.551961
Rsn62_27 sn62_27 sn63_27 11.551961
Rsp62_28 sp62_28 sp63_28 11.551961
Rsn62_28 sn62_28 sn63_28 11.551961
Rsp62_29 sp62_29 sp63_29 11.551961
Rsn62_29 sn62_29 sn63_29 11.551961
Rsp62_30 sp62_30 sp63_30 11.551961
Rsn62_30 sn62_30 sn63_30 11.551961
Rsp62_31 sp62_31 sp63_31 11.551961
Rsn62_31 sn62_31 sn63_31 11.551961
Rsp62_32 sp62_32 sp63_32 11.551961
Rsn62_32 sn62_32 sn63_32 11.551961
Rsp62_33 sp62_33 sp63_33 11.551961
Rsn62_33 sn62_33 sn63_33 11.551961
Rsp62_34 sp62_34 sp63_34 11.551961
Rsn62_34 sn62_34 sn63_34 11.551961
Rsp62_35 sp62_35 sp63_35 11.551961
Rsn62_35 sn62_35 sn63_35 11.551961
Rsp62_36 sp62_36 sp63_36 11.551961
Rsn62_36 sn62_36 sn63_36 11.551961
Rsp62_37 sp62_37 sp63_37 11.551961
Rsn62_37 sn62_37 sn63_37 11.551961
Rsp62_38 sp62_38 sp63_38 11.551961
Rsn62_38 sn62_38 sn63_38 11.551961
Rsp62_39 sp62_39 sp63_39 11.551961
Rsn62_39 sn62_39 sn63_39 11.551961
Rsp62_40 sp62_40 sp63_40 11.551961
Rsn62_40 sn62_40 sn63_40 11.551961
Rsp62_41 sp62_41 sp63_41 11.551961
Rsn62_41 sn62_41 sn63_41 11.551961
Rsp62_42 sp62_42 sp63_42 11.551961
Rsn62_42 sn62_42 sn63_42 11.551961
Rsp62_43 sp62_43 sp63_43 11.551961
Rsn62_43 sn62_43 sn63_43 11.551961
Rsp62_44 sp62_44 sp63_44 11.551961
Rsn62_44 sn62_44 sn63_44 11.551961
Rsp62_45 sp62_45 sp63_45 11.551961
Rsn62_45 sn62_45 sn63_45 11.551961
Rsp62_46 sp62_46 sp63_46 11.551961
Rsn62_46 sn62_46 sn63_46 11.551961
Rsp62_47 sp62_47 sp63_47 11.551961
Rsn62_47 sn62_47 sn63_47 11.551961
Rsp62_48 sp62_48 sp63_48 11.551961
Rsn62_48 sn62_48 sn63_48 11.551961
Rsp62_49 sp62_49 sp63_49 11.551961
Rsn62_49 sn62_49 sn63_49 11.551961
Rsp62_50 sp62_50 sp63_50 11.551961
Rsn62_50 sn62_50 sn63_50 11.551961
Rsp62_51 sp62_51 sp63_51 11.551961
Rsn62_51 sn62_51 sn63_51 11.551961
Rsp62_52 sp62_52 sp63_52 11.551961
Rsn62_52 sn62_52 sn63_52 11.551961
Rsp62_53 sp62_53 sp63_53 11.551961
Rsn62_53 sn62_53 sn63_53 11.551961
Rsp62_54 sp62_54 sp63_54 11.551961
Rsn62_54 sn62_54 sn63_54 11.551961
Rsp62_55 sp62_55 sp63_55 11.551961
Rsn62_55 sn62_55 sn63_55 11.551961
Rsp62_56 sp62_56 sp63_56 11.551961
Rsn62_56 sn62_56 sn63_56 11.551961
Rsp62_57 sp62_57 sp63_57 11.551961
Rsn62_57 sn62_57 sn63_57 11.551961
Rsp62_58 sp62_58 sp63_58 11.551961
Rsn62_58 sn62_58 sn63_58 11.551961
Rsp62_59 sp62_59 sp63_59 11.551961
Rsn62_59 sn62_59 sn63_59 11.551961
Rsp62_60 sp62_60 sp63_60 11.551961
Rsn62_60 sn62_60 sn63_60 11.551961
Rsp62_61 sp62_61 sp63_61 11.551961
Rsn62_61 sn62_61 sn63_61 11.551961
Rsp62_62 sp62_62 sp63_62 11.551961
Rsn62_62 sn62_62 sn63_62 11.551961
Rsp62_63 sp62_63 sp63_63 11.551961
Rsn62_63 sn62_63 sn63_63 11.551961
Rsp62_64 sp62_64 sp63_64 11.551961
Rsn62_64 sn62_64 sn63_64 11.551961
Rsp62_65 sp62_65 sp63_65 11.551961
Rsn62_65 sn62_65 sn63_65 11.551961
Rsp62_66 sp62_66 sp63_66 11.551961
Rsn62_66 sn62_66 sn63_66 11.551961
Rsp62_67 sp62_67 sp63_67 11.551961
Rsn62_67 sn62_67 sn63_67 11.551961
Rsp62_68 sp62_68 sp63_68 11.551961
Rsn62_68 sn62_68 sn63_68 11.551961
Rsp62_69 sp62_69 sp63_69 11.551961
Rsn62_69 sn62_69 sn63_69 11.551961
Rsp62_70 sp62_70 sp63_70 11.551961
Rsn62_70 sn62_70 sn63_70 11.551961
Rsp62_71 sp62_71 sp63_71 11.551961
Rsn62_71 sn62_71 sn63_71 11.551961
Rsp62_72 sp62_72 sp63_72 11.551961
Rsn62_72 sn62_72 sn63_72 11.551961
Rsp62_73 sp62_73 sp63_73 11.551961
Rsn62_73 sn62_73 sn63_73 11.551961
Rsp62_74 sp62_74 sp63_74 11.551961
Rsn62_74 sn62_74 sn63_74 11.551961
Rsp62_75 sp62_75 sp63_75 11.551961
Rsn62_75 sn62_75 sn63_75 11.551961
Rsp62_76 sp62_76 sp63_76 11.551961
Rsn62_76 sn62_76 sn63_76 11.551961
Rsp62_77 sp62_77 sp63_77 11.551961
Rsn62_77 sn62_77 sn63_77 11.551961
Rsp62_78 sp62_78 sp63_78 11.551961
Rsn62_78 sn62_78 sn63_78 11.551961
Rsp62_79 sp62_79 sp63_79 11.551961
Rsn62_79 sn62_79 sn63_79 11.551961
Rsp62_80 sp62_80 sp63_80 11.551961
Rsn62_80 sn62_80 sn63_80 11.551961
Rsp62_81 sp62_81 sp63_81 11.551961
Rsn62_81 sn62_81 sn63_81 11.551961
Rsp62_82 sp62_82 sp63_82 11.551961
Rsn62_82 sn62_82 sn63_82 11.551961
Rsp62_83 sp62_83 sp63_83 11.551961
Rsn62_83 sn62_83 sn63_83 11.551961
Rsp62_84 sp62_84 sp63_84 11.551961
Rsn62_84 sn62_84 sn63_84 11.551961
Rsp63_1 sp63_1 sp64_1 11.551961
Rsn63_1 sn63_1 sn64_1 11.551961
Rsp63_2 sp63_2 sp64_2 11.551961
Rsn63_2 sn63_2 sn64_2 11.551961
Rsp63_3 sp63_3 sp64_3 11.551961
Rsn63_3 sn63_3 sn64_3 11.551961
Rsp63_4 sp63_4 sp64_4 11.551961
Rsn63_4 sn63_4 sn64_4 11.551961
Rsp63_5 sp63_5 sp64_5 11.551961
Rsn63_5 sn63_5 sn64_5 11.551961
Rsp63_6 sp63_6 sp64_6 11.551961
Rsn63_6 sn63_6 sn64_6 11.551961
Rsp63_7 sp63_7 sp64_7 11.551961
Rsn63_7 sn63_7 sn64_7 11.551961
Rsp63_8 sp63_8 sp64_8 11.551961
Rsn63_8 sn63_8 sn64_8 11.551961
Rsp63_9 sp63_9 sp64_9 11.551961
Rsn63_9 sn63_9 sn64_9 11.551961
Rsp63_10 sp63_10 sp64_10 11.551961
Rsn63_10 sn63_10 sn64_10 11.551961
Rsp63_11 sp63_11 sp64_11 11.551961
Rsn63_11 sn63_11 sn64_11 11.551961
Rsp63_12 sp63_12 sp64_12 11.551961
Rsn63_12 sn63_12 sn64_12 11.551961
Rsp63_13 sp63_13 sp64_13 11.551961
Rsn63_13 sn63_13 sn64_13 11.551961
Rsp63_14 sp63_14 sp64_14 11.551961
Rsn63_14 sn63_14 sn64_14 11.551961
Rsp63_15 sp63_15 sp64_15 11.551961
Rsn63_15 sn63_15 sn64_15 11.551961
Rsp63_16 sp63_16 sp64_16 11.551961
Rsn63_16 sn63_16 sn64_16 11.551961
Rsp63_17 sp63_17 sp64_17 11.551961
Rsn63_17 sn63_17 sn64_17 11.551961
Rsp63_18 sp63_18 sp64_18 11.551961
Rsn63_18 sn63_18 sn64_18 11.551961
Rsp63_19 sp63_19 sp64_19 11.551961
Rsn63_19 sn63_19 sn64_19 11.551961
Rsp63_20 sp63_20 sp64_20 11.551961
Rsn63_20 sn63_20 sn64_20 11.551961
Rsp63_21 sp63_21 sp64_21 11.551961
Rsn63_21 sn63_21 sn64_21 11.551961
Rsp63_22 sp63_22 sp64_22 11.551961
Rsn63_22 sn63_22 sn64_22 11.551961
Rsp63_23 sp63_23 sp64_23 11.551961
Rsn63_23 sn63_23 sn64_23 11.551961
Rsp63_24 sp63_24 sp64_24 11.551961
Rsn63_24 sn63_24 sn64_24 11.551961
Rsp63_25 sp63_25 sp64_25 11.551961
Rsn63_25 sn63_25 sn64_25 11.551961
Rsp63_26 sp63_26 sp64_26 11.551961
Rsn63_26 sn63_26 sn64_26 11.551961
Rsp63_27 sp63_27 sp64_27 11.551961
Rsn63_27 sn63_27 sn64_27 11.551961
Rsp63_28 sp63_28 sp64_28 11.551961
Rsn63_28 sn63_28 sn64_28 11.551961
Rsp63_29 sp63_29 sp64_29 11.551961
Rsn63_29 sn63_29 sn64_29 11.551961
Rsp63_30 sp63_30 sp64_30 11.551961
Rsn63_30 sn63_30 sn64_30 11.551961
Rsp63_31 sp63_31 sp64_31 11.551961
Rsn63_31 sn63_31 sn64_31 11.551961
Rsp63_32 sp63_32 sp64_32 11.551961
Rsn63_32 sn63_32 sn64_32 11.551961
Rsp63_33 sp63_33 sp64_33 11.551961
Rsn63_33 sn63_33 sn64_33 11.551961
Rsp63_34 sp63_34 sp64_34 11.551961
Rsn63_34 sn63_34 sn64_34 11.551961
Rsp63_35 sp63_35 sp64_35 11.551961
Rsn63_35 sn63_35 sn64_35 11.551961
Rsp63_36 sp63_36 sp64_36 11.551961
Rsn63_36 sn63_36 sn64_36 11.551961
Rsp63_37 sp63_37 sp64_37 11.551961
Rsn63_37 sn63_37 sn64_37 11.551961
Rsp63_38 sp63_38 sp64_38 11.551961
Rsn63_38 sn63_38 sn64_38 11.551961
Rsp63_39 sp63_39 sp64_39 11.551961
Rsn63_39 sn63_39 sn64_39 11.551961
Rsp63_40 sp63_40 sp64_40 11.551961
Rsn63_40 sn63_40 sn64_40 11.551961
Rsp63_41 sp63_41 sp64_41 11.551961
Rsn63_41 sn63_41 sn64_41 11.551961
Rsp63_42 sp63_42 sp64_42 11.551961
Rsn63_42 sn63_42 sn64_42 11.551961
Rsp63_43 sp63_43 sp64_43 11.551961
Rsn63_43 sn63_43 sn64_43 11.551961
Rsp63_44 sp63_44 sp64_44 11.551961
Rsn63_44 sn63_44 sn64_44 11.551961
Rsp63_45 sp63_45 sp64_45 11.551961
Rsn63_45 sn63_45 sn64_45 11.551961
Rsp63_46 sp63_46 sp64_46 11.551961
Rsn63_46 sn63_46 sn64_46 11.551961
Rsp63_47 sp63_47 sp64_47 11.551961
Rsn63_47 sn63_47 sn64_47 11.551961
Rsp63_48 sp63_48 sp64_48 11.551961
Rsn63_48 sn63_48 sn64_48 11.551961
Rsp63_49 sp63_49 sp64_49 11.551961
Rsn63_49 sn63_49 sn64_49 11.551961
Rsp63_50 sp63_50 sp64_50 11.551961
Rsn63_50 sn63_50 sn64_50 11.551961
Rsp63_51 sp63_51 sp64_51 11.551961
Rsn63_51 sn63_51 sn64_51 11.551961
Rsp63_52 sp63_52 sp64_52 11.551961
Rsn63_52 sn63_52 sn64_52 11.551961
Rsp63_53 sp63_53 sp64_53 11.551961
Rsn63_53 sn63_53 sn64_53 11.551961
Rsp63_54 sp63_54 sp64_54 11.551961
Rsn63_54 sn63_54 sn64_54 11.551961
Rsp63_55 sp63_55 sp64_55 11.551961
Rsn63_55 sn63_55 sn64_55 11.551961
Rsp63_56 sp63_56 sp64_56 11.551961
Rsn63_56 sn63_56 sn64_56 11.551961
Rsp63_57 sp63_57 sp64_57 11.551961
Rsn63_57 sn63_57 sn64_57 11.551961
Rsp63_58 sp63_58 sp64_58 11.551961
Rsn63_58 sn63_58 sn64_58 11.551961
Rsp63_59 sp63_59 sp64_59 11.551961
Rsn63_59 sn63_59 sn64_59 11.551961
Rsp63_60 sp63_60 sp64_60 11.551961
Rsn63_60 sn63_60 sn64_60 11.551961
Rsp63_61 sp63_61 sp64_61 11.551961
Rsn63_61 sn63_61 sn64_61 11.551961
Rsp63_62 sp63_62 sp64_62 11.551961
Rsn63_62 sn63_62 sn64_62 11.551961
Rsp63_63 sp63_63 sp64_63 11.551961
Rsn63_63 sn63_63 sn64_63 11.551961
Rsp63_64 sp63_64 sp64_64 11.551961
Rsn63_64 sn63_64 sn64_64 11.551961
Rsp63_65 sp63_65 sp64_65 11.551961
Rsn63_65 sn63_65 sn64_65 11.551961
Rsp63_66 sp63_66 sp64_66 11.551961
Rsn63_66 sn63_66 sn64_66 11.551961
Rsp63_67 sp63_67 sp64_67 11.551961
Rsn63_67 sn63_67 sn64_67 11.551961
Rsp63_68 sp63_68 sp64_68 11.551961
Rsn63_68 sn63_68 sn64_68 11.551961
Rsp63_69 sp63_69 sp64_69 11.551961
Rsn63_69 sn63_69 sn64_69 11.551961
Rsp63_70 sp63_70 sp64_70 11.551961
Rsn63_70 sn63_70 sn64_70 11.551961
Rsp63_71 sp63_71 sp64_71 11.551961
Rsn63_71 sn63_71 sn64_71 11.551961
Rsp63_72 sp63_72 sp64_72 11.551961
Rsn63_72 sn63_72 sn64_72 11.551961
Rsp63_73 sp63_73 sp64_73 11.551961
Rsn63_73 sn63_73 sn64_73 11.551961
Rsp63_74 sp63_74 sp64_74 11.551961
Rsn63_74 sn63_74 sn64_74 11.551961
Rsp63_75 sp63_75 sp64_75 11.551961
Rsn63_75 sn63_75 sn64_75 11.551961
Rsp63_76 sp63_76 sp64_76 11.551961
Rsn63_76 sn63_76 sn64_76 11.551961
Rsp63_77 sp63_77 sp64_77 11.551961
Rsn63_77 sn63_77 sn64_77 11.551961
Rsp63_78 sp63_78 sp64_78 11.551961
Rsn63_78 sn63_78 sn64_78 11.551961
Rsp63_79 sp63_79 sp64_79 11.551961
Rsn63_79 sn63_79 sn64_79 11.551961
Rsp63_80 sp63_80 sp64_80 11.551961
Rsn63_80 sn63_80 sn64_80 11.551961
Rsp63_81 sp63_81 sp64_81 11.551961
Rsn63_81 sn63_81 sn64_81 11.551961
Rsp63_82 sp63_82 sp64_82 11.551961
Rsn63_82 sn63_82 sn64_82 11.551961
Rsp63_83 sp63_83 sp64_83 11.551961
Rsn63_83 sn63_83 sn64_83 11.551961
Rsp63_84 sp63_84 sp64_84 11.551961
Rsn63_84 sn63_84 sn64_84 11.551961
Rsp64_1 sp64_1 sp65_1 11.551961
Rsn64_1 sn64_1 sn65_1 11.551961
Rsp64_2 sp64_2 sp65_2 11.551961
Rsn64_2 sn64_2 sn65_2 11.551961
Rsp64_3 sp64_3 sp65_3 11.551961
Rsn64_3 sn64_3 sn65_3 11.551961
Rsp64_4 sp64_4 sp65_4 11.551961
Rsn64_4 sn64_4 sn65_4 11.551961
Rsp64_5 sp64_5 sp65_5 11.551961
Rsn64_5 sn64_5 sn65_5 11.551961
Rsp64_6 sp64_6 sp65_6 11.551961
Rsn64_6 sn64_6 sn65_6 11.551961
Rsp64_7 sp64_7 sp65_7 11.551961
Rsn64_7 sn64_7 sn65_7 11.551961
Rsp64_8 sp64_8 sp65_8 11.551961
Rsn64_8 sn64_8 sn65_8 11.551961
Rsp64_9 sp64_9 sp65_9 11.551961
Rsn64_9 sn64_9 sn65_9 11.551961
Rsp64_10 sp64_10 sp65_10 11.551961
Rsn64_10 sn64_10 sn65_10 11.551961
Rsp64_11 sp64_11 sp65_11 11.551961
Rsn64_11 sn64_11 sn65_11 11.551961
Rsp64_12 sp64_12 sp65_12 11.551961
Rsn64_12 sn64_12 sn65_12 11.551961
Rsp64_13 sp64_13 sp65_13 11.551961
Rsn64_13 sn64_13 sn65_13 11.551961
Rsp64_14 sp64_14 sp65_14 11.551961
Rsn64_14 sn64_14 sn65_14 11.551961
Rsp64_15 sp64_15 sp65_15 11.551961
Rsn64_15 sn64_15 sn65_15 11.551961
Rsp64_16 sp64_16 sp65_16 11.551961
Rsn64_16 sn64_16 sn65_16 11.551961
Rsp64_17 sp64_17 sp65_17 11.551961
Rsn64_17 sn64_17 sn65_17 11.551961
Rsp64_18 sp64_18 sp65_18 11.551961
Rsn64_18 sn64_18 sn65_18 11.551961
Rsp64_19 sp64_19 sp65_19 11.551961
Rsn64_19 sn64_19 sn65_19 11.551961
Rsp64_20 sp64_20 sp65_20 11.551961
Rsn64_20 sn64_20 sn65_20 11.551961
Rsp64_21 sp64_21 sp65_21 11.551961
Rsn64_21 sn64_21 sn65_21 11.551961
Rsp64_22 sp64_22 sp65_22 11.551961
Rsn64_22 sn64_22 sn65_22 11.551961
Rsp64_23 sp64_23 sp65_23 11.551961
Rsn64_23 sn64_23 sn65_23 11.551961
Rsp64_24 sp64_24 sp65_24 11.551961
Rsn64_24 sn64_24 sn65_24 11.551961
Rsp64_25 sp64_25 sp65_25 11.551961
Rsn64_25 sn64_25 sn65_25 11.551961
Rsp64_26 sp64_26 sp65_26 11.551961
Rsn64_26 sn64_26 sn65_26 11.551961
Rsp64_27 sp64_27 sp65_27 11.551961
Rsn64_27 sn64_27 sn65_27 11.551961
Rsp64_28 sp64_28 sp65_28 11.551961
Rsn64_28 sn64_28 sn65_28 11.551961
Rsp64_29 sp64_29 sp65_29 11.551961
Rsn64_29 sn64_29 sn65_29 11.551961
Rsp64_30 sp64_30 sp65_30 11.551961
Rsn64_30 sn64_30 sn65_30 11.551961
Rsp64_31 sp64_31 sp65_31 11.551961
Rsn64_31 sn64_31 sn65_31 11.551961
Rsp64_32 sp64_32 sp65_32 11.551961
Rsn64_32 sn64_32 sn65_32 11.551961
Rsp64_33 sp64_33 sp65_33 11.551961
Rsn64_33 sn64_33 sn65_33 11.551961
Rsp64_34 sp64_34 sp65_34 11.551961
Rsn64_34 sn64_34 sn65_34 11.551961
Rsp64_35 sp64_35 sp65_35 11.551961
Rsn64_35 sn64_35 sn65_35 11.551961
Rsp64_36 sp64_36 sp65_36 11.551961
Rsn64_36 sn64_36 sn65_36 11.551961
Rsp64_37 sp64_37 sp65_37 11.551961
Rsn64_37 sn64_37 sn65_37 11.551961
Rsp64_38 sp64_38 sp65_38 11.551961
Rsn64_38 sn64_38 sn65_38 11.551961
Rsp64_39 sp64_39 sp65_39 11.551961
Rsn64_39 sn64_39 sn65_39 11.551961
Rsp64_40 sp64_40 sp65_40 11.551961
Rsn64_40 sn64_40 sn65_40 11.551961
Rsp64_41 sp64_41 sp65_41 11.551961
Rsn64_41 sn64_41 sn65_41 11.551961
Rsp64_42 sp64_42 sp65_42 11.551961
Rsn64_42 sn64_42 sn65_42 11.551961
Rsp64_43 sp64_43 sp65_43 11.551961
Rsn64_43 sn64_43 sn65_43 11.551961
Rsp64_44 sp64_44 sp65_44 11.551961
Rsn64_44 sn64_44 sn65_44 11.551961
Rsp64_45 sp64_45 sp65_45 11.551961
Rsn64_45 sn64_45 sn65_45 11.551961
Rsp64_46 sp64_46 sp65_46 11.551961
Rsn64_46 sn64_46 sn65_46 11.551961
Rsp64_47 sp64_47 sp65_47 11.551961
Rsn64_47 sn64_47 sn65_47 11.551961
Rsp64_48 sp64_48 sp65_48 11.551961
Rsn64_48 sn64_48 sn65_48 11.551961
Rsp64_49 sp64_49 sp65_49 11.551961
Rsn64_49 sn64_49 sn65_49 11.551961
Rsp64_50 sp64_50 sp65_50 11.551961
Rsn64_50 sn64_50 sn65_50 11.551961
Rsp64_51 sp64_51 sp65_51 11.551961
Rsn64_51 sn64_51 sn65_51 11.551961
Rsp64_52 sp64_52 sp65_52 11.551961
Rsn64_52 sn64_52 sn65_52 11.551961
Rsp64_53 sp64_53 sp65_53 11.551961
Rsn64_53 sn64_53 sn65_53 11.551961
Rsp64_54 sp64_54 sp65_54 11.551961
Rsn64_54 sn64_54 sn65_54 11.551961
Rsp64_55 sp64_55 sp65_55 11.551961
Rsn64_55 sn64_55 sn65_55 11.551961
Rsp64_56 sp64_56 sp65_56 11.551961
Rsn64_56 sn64_56 sn65_56 11.551961
Rsp64_57 sp64_57 sp65_57 11.551961
Rsn64_57 sn64_57 sn65_57 11.551961
Rsp64_58 sp64_58 sp65_58 11.551961
Rsn64_58 sn64_58 sn65_58 11.551961
Rsp64_59 sp64_59 sp65_59 11.551961
Rsn64_59 sn64_59 sn65_59 11.551961
Rsp64_60 sp64_60 sp65_60 11.551961
Rsn64_60 sn64_60 sn65_60 11.551961
Rsp64_61 sp64_61 sp65_61 11.551961
Rsn64_61 sn64_61 sn65_61 11.551961
Rsp64_62 sp64_62 sp65_62 11.551961
Rsn64_62 sn64_62 sn65_62 11.551961
Rsp64_63 sp64_63 sp65_63 11.551961
Rsn64_63 sn64_63 sn65_63 11.551961
Rsp64_64 sp64_64 sp65_64 11.551961
Rsn64_64 sn64_64 sn65_64 11.551961
Rsp64_65 sp64_65 sp65_65 11.551961
Rsn64_65 sn64_65 sn65_65 11.551961
Rsp64_66 sp64_66 sp65_66 11.551961
Rsn64_66 sn64_66 sn65_66 11.551961
Rsp64_67 sp64_67 sp65_67 11.551961
Rsn64_67 sn64_67 sn65_67 11.551961
Rsp64_68 sp64_68 sp65_68 11.551961
Rsn64_68 sn64_68 sn65_68 11.551961
Rsp64_69 sp64_69 sp65_69 11.551961
Rsn64_69 sn64_69 sn65_69 11.551961
Rsp64_70 sp64_70 sp65_70 11.551961
Rsn64_70 sn64_70 sn65_70 11.551961
Rsp64_71 sp64_71 sp65_71 11.551961
Rsn64_71 sn64_71 sn65_71 11.551961
Rsp64_72 sp64_72 sp65_72 11.551961
Rsn64_72 sn64_72 sn65_72 11.551961
Rsp64_73 sp64_73 sp65_73 11.551961
Rsn64_73 sn64_73 sn65_73 11.551961
Rsp64_74 sp64_74 sp65_74 11.551961
Rsn64_74 sn64_74 sn65_74 11.551961
Rsp64_75 sp64_75 sp65_75 11.551961
Rsn64_75 sn64_75 sn65_75 11.551961
Rsp64_76 sp64_76 sp65_76 11.551961
Rsn64_76 sn64_76 sn65_76 11.551961
Rsp64_77 sp64_77 sp65_77 11.551961
Rsn64_77 sn64_77 sn65_77 11.551961
Rsp64_78 sp64_78 sp65_78 11.551961
Rsn64_78 sn64_78 sn65_78 11.551961
Rsp64_79 sp64_79 sp65_79 11.551961
Rsn64_79 sn64_79 sn65_79 11.551961
Rsp64_80 sp64_80 sp65_80 11.551961
Rsn64_80 sn64_80 sn65_80 11.551961
Rsp64_81 sp64_81 sp65_81 11.551961
Rsn64_81 sn64_81 sn65_81 11.551961
Rsp64_82 sp64_82 sp65_82 11.551961
Rsn64_82 sn64_82 sn65_82 11.551961
Rsp64_83 sp64_83 sp65_83 11.551961
Rsn64_83 sn64_83 sn65_83 11.551961
Rsp64_84 sp64_84 sp65_84 11.551961
Rsn64_84 sn64_84 sn65_84 11.551961
Rsp65_1 sp65_1 sp66_1 11.551961
Rsn65_1 sn65_1 sn66_1 11.551961
Rsp65_2 sp65_2 sp66_2 11.551961
Rsn65_2 sn65_2 sn66_2 11.551961
Rsp65_3 sp65_3 sp66_3 11.551961
Rsn65_3 sn65_3 sn66_3 11.551961
Rsp65_4 sp65_4 sp66_4 11.551961
Rsn65_4 sn65_4 sn66_4 11.551961
Rsp65_5 sp65_5 sp66_5 11.551961
Rsn65_5 sn65_5 sn66_5 11.551961
Rsp65_6 sp65_6 sp66_6 11.551961
Rsn65_6 sn65_6 sn66_6 11.551961
Rsp65_7 sp65_7 sp66_7 11.551961
Rsn65_7 sn65_7 sn66_7 11.551961
Rsp65_8 sp65_8 sp66_8 11.551961
Rsn65_8 sn65_8 sn66_8 11.551961
Rsp65_9 sp65_9 sp66_9 11.551961
Rsn65_9 sn65_9 sn66_9 11.551961
Rsp65_10 sp65_10 sp66_10 11.551961
Rsn65_10 sn65_10 sn66_10 11.551961
Rsp65_11 sp65_11 sp66_11 11.551961
Rsn65_11 sn65_11 sn66_11 11.551961
Rsp65_12 sp65_12 sp66_12 11.551961
Rsn65_12 sn65_12 sn66_12 11.551961
Rsp65_13 sp65_13 sp66_13 11.551961
Rsn65_13 sn65_13 sn66_13 11.551961
Rsp65_14 sp65_14 sp66_14 11.551961
Rsn65_14 sn65_14 sn66_14 11.551961
Rsp65_15 sp65_15 sp66_15 11.551961
Rsn65_15 sn65_15 sn66_15 11.551961
Rsp65_16 sp65_16 sp66_16 11.551961
Rsn65_16 sn65_16 sn66_16 11.551961
Rsp65_17 sp65_17 sp66_17 11.551961
Rsn65_17 sn65_17 sn66_17 11.551961
Rsp65_18 sp65_18 sp66_18 11.551961
Rsn65_18 sn65_18 sn66_18 11.551961
Rsp65_19 sp65_19 sp66_19 11.551961
Rsn65_19 sn65_19 sn66_19 11.551961
Rsp65_20 sp65_20 sp66_20 11.551961
Rsn65_20 sn65_20 sn66_20 11.551961
Rsp65_21 sp65_21 sp66_21 11.551961
Rsn65_21 sn65_21 sn66_21 11.551961
Rsp65_22 sp65_22 sp66_22 11.551961
Rsn65_22 sn65_22 sn66_22 11.551961
Rsp65_23 sp65_23 sp66_23 11.551961
Rsn65_23 sn65_23 sn66_23 11.551961
Rsp65_24 sp65_24 sp66_24 11.551961
Rsn65_24 sn65_24 sn66_24 11.551961
Rsp65_25 sp65_25 sp66_25 11.551961
Rsn65_25 sn65_25 sn66_25 11.551961
Rsp65_26 sp65_26 sp66_26 11.551961
Rsn65_26 sn65_26 sn66_26 11.551961
Rsp65_27 sp65_27 sp66_27 11.551961
Rsn65_27 sn65_27 sn66_27 11.551961
Rsp65_28 sp65_28 sp66_28 11.551961
Rsn65_28 sn65_28 sn66_28 11.551961
Rsp65_29 sp65_29 sp66_29 11.551961
Rsn65_29 sn65_29 sn66_29 11.551961
Rsp65_30 sp65_30 sp66_30 11.551961
Rsn65_30 sn65_30 sn66_30 11.551961
Rsp65_31 sp65_31 sp66_31 11.551961
Rsn65_31 sn65_31 sn66_31 11.551961
Rsp65_32 sp65_32 sp66_32 11.551961
Rsn65_32 sn65_32 sn66_32 11.551961
Rsp65_33 sp65_33 sp66_33 11.551961
Rsn65_33 sn65_33 sn66_33 11.551961
Rsp65_34 sp65_34 sp66_34 11.551961
Rsn65_34 sn65_34 sn66_34 11.551961
Rsp65_35 sp65_35 sp66_35 11.551961
Rsn65_35 sn65_35 sn66_35 11.551961
Rsp65_36 sp65_36 sp66_36 11.551961
Rsn65_36 sn65_36 sn66_36 11.551961
Rsp65_37 sp65_37 sp66_37 11.551961
Rsn65_37 sn65_37 sn66_37 11.551961
Rsp65_38 sp65_38 sp66_38 11.551961
Rsn65_38 sn65_38 sn66_38 11.551961
Rsp65_39 sp65_39 sp66_39 11.551961
Rsn65_39 sn65_39 sn66_39 11.551961
Rsp65_40 sp65_40 sp66_40 11.551961
Rsn65_40 sn65_40 sn66_40 11.551961
Rsp65_41 sp65_41 sp66_41 11.551961
Rsn65_41 sn65_41 sn66_41 11.551961
Rsp65_42 sp65_42 sp66_42 11.551961
Rsn65_42 sn65_42 sn66_42 11.551961
Rsp65_43 sp65_43 sp66_43 11.551961
Rsn65_43 sn65_43 sn66_43 11.551961
Rsp65_44 sp65_44 sp66_44 11.551961
Rsn65_44 sn65_44 sn66_44 11.551961
Rsp65_45 sp65_45 sp66_45 11.551961
Rsn65_45 sn65_45 sn66_45 11.551961
Rsp65_46 sp65_46 sp66_46 11.551961
Rsn65_46 sn65_46 sn66_46 11.551961
Rsp65_47 sp65_47 sp66_47 11.551961
Rsn65_47 sn65_47 sn66_47 11.551961
Rsp65_48 sp65_48 sp66_48 11.551961
Rsn65_48 sn65_48 sn66_48 11.551961
Rsp65_49 sp65_49 sp66_49 11.551961
Rsn65_49 sn65_49 sn66_49 11.551961
Rsp65_50 sp65_50 sp66_50 11.551961
Rsn65_50 sn65_50 sn66_50 11.551961
Rsp65_51 sp65_51 sp66_51 11.551961
Rsn65_51 sn65_51 sn66_51 11.551961
Rsp65_52 sp65_52 sp66_52 11.551961
Rsn65_52 sn65_52 sn66_52 11.551961
Rsp65_53 sp65_53 sp66_53 11.551961
Rsn65_53 sn65_53 sn66_53 11.551961
Rsp65_54 sp65_54 sp66_54 11.551961
Rsn65_54 sn65_54 sn66_54 11.551961
Rsp65_55 sp65_55 sp66_55 11.551961
Rsn65_55 sn65_55 sn66_55 11.551961
Rsp65_56 sp65_56 sp66_56 11.551961
Rsn65_56 sn65_56 sn66_56 11.551961
Rsp65_57 sp65_57 sp66_57 11.551961
Rsn65_57 sn65_57 sn66_57 11.551961
Rsp65_58 sp65_58 sp66_58 11.551961
Rsn65_58 sn65_58 sn66_58 11.551961
Rsp65_59 sp65_59 sp66_59 11.551961
Rsn65_59 sn65_59 sn66_59 11.551961
Rsp65_60 sp65_60 sp66_60 11.551961
Rsn65_60 sn65_60 sn66_60 11.551961
Rsp65_61 sp65_61 sp66_61 11.551961
Rsn65_61 sn65_61 sn66_61 11.551961
Rsp65_62 sp65_62 sp66_62 11.551961
Rsn65_62 sn65_62 sn66_62 11.551961
Rsp65_63 sp65_63 sp66_63 11.551961
Rsn65_63 sn65_63 sn66_63 11.551961
Rsp65_64 sp65_64 sp66_64 11.551961
Rsn65_64 sn65_64 sn66_64 11.551961
Rsp65_65 sp65_65 sp66_65 11.551961
Rsn65_65 sn65_65 sn66_65 11.551961
Rsp65_66 sp65_66 sp66_66 11.551961
Rsn65_66 sn65_66 sn66_66 11.551961
Rsp65_67 sp65_67 sp66_67 11.551961
Rsn65_67 sn65_67 sn66_67 11.551961
Rsp65_68 sp65_68 sp66_68 11.551961
Rsn65_68 sn65_68 sn66_68 11.551961
Rsp65_69 sp65_69 sp66_69 11.551961
Rsn65_69 sn65_69 sn66_69 11.551961
Rsp65_70 sp65_70 sp66_70 11.551961
Rsn65_70 sn65_70 sn66_70 11.551961
Rsp65_71 sp65_71 sp66_71 11.551961
Rsn65_71 sn65_71 sn66_71 11.551961
Rsp65_72 sp65_72 sp66_72 11.551961
Rsn65_72 sn65_72 sn66_72 11.551961
Rsp65_73 sp65_73 sp66_73 11.551961
Rsn65_73 sn65_73 sn66_73 11.551961
Rsp65_74 sp65_74 sp66_74 11.551961
Rsn65_74 sn65_74 sn66_74 11.551961
Rsp65_75 sp65_75 sp66_75 11.551961
Rsn65_75 sn65_75 sn66_75 11.551961
Rsp65_76 sp65_76 sp66_76 11.551961
Rsn65_76 sn65_76 sn66_76 11.551961
Rsp65_77 sp65_77 sp66_77 11.551961
Rsn65_77 sn65_77 sn66_77 11.551961
Rsp65_78 sp65_78 sp66_78 11.551961
Rsn65_78 sn65_78 sn66_78 11.551961
Rsp65_79 sp65_79 sp66_79 11.551961
Rsn65_79 sn65_79 sn66_79 11.551961
Rsp65_80 sp65_80 sp66_80 11.551961
Rsn65_80 sn65_80 sn66_80 11.551961
Rsp65_81 sp65_81 sp66_81 11.551961
Rsn65_81 sn65_81 sn66_81 11.551961
Rsp65_82 sp65_82 sp66_82 11.551961
Rsn65_82 sn65_82 sn66_82 11.551961
Rsp65_83 sp65_83 sp66_83 11.551961
Rsn65_83 sn65_83 sn66_83 11.551961
Rsp65_84 sp65_84 sp66_84 11.551961
Rsn65_84 sn65_84 sn66_84 11.551961
Rsp66_1 sp66_1 sp67_1 11.551961
Rsn66_1 sn66_1 sn67_1 11.551961
Rsp66_2 sp66_2 sp67_2 11.551961
Rsn66_2 sn66_2 sn67_2 11.551961
Rsp66_3 sp66_3 sp67_3 11.551961
Rsn66_3 sn66_3 sn67_3 11.551961
Rsp66_4 sp66_4 sp67_4 11.551961
Rsn66_4 sn66_4 sn67_4 11.551961
Rsp66_5 sp66_5 sp67_5 11.551961
Rsn66_5 sn66_5 sn67_5 11.551961
Rsp66_6 sp66_6 sp67_6 11.551961
Rsn66_6 sn66_6 sn67_6 11.551961
Rsp66_7 sp66_7 sp67_7 11.551961
Rsn66_7 sn66_7 sn67_7 11.551961
Rsp66_8 sp66_8 sp67_8 11.551961
Rsn66_8 sn66_8 sn67_8 11.551961
Rsp66_9 sp66_9 sp67_9 11.551961
Rsn66_9 sn66_9 sn67_9 11.551961
Rsp66_10 sp66_10 sp67_10 11.551961
Rsn66_10 sn66_10 sn67_10 11.551961
Rsp66_11 sp66_11 sp67_11 11.551961
Rsn66_11 sn66_11 sn67_11 11.551961
Rsp66_12 sp66_12 sp67_12 11.551961
Rsn66_12 sn66_12 sn67_12 11.551961
Rsp66_13 sp66_13 sp67_13 11.551961
Rsn66_13 sn66_13 sn67_13 11.551961
Rsp66_14 sp66_14 sp67_14 11.551961
Rsn66_14 sn66_14 sn67_14 11.551961
Rsp66_15 sp66_15 sp67_15 11.551961
Rsn66_15 sn66_15 sn67_15 11.551961
Rsp66_16 sp66_16 sp67_16 11.551961
Rsn66_16 sn66_16 sn67_16 11.551961
Rsp66_17 sp66_17 sp67_17 11.551961
Rsn66_17 sn66_17 sn67_17 11.551961
Rsp66_18 sp66_18 sp67_18 11.551961
Rsn66_18 sn66_18 sn67_18 11.551961
Rsp66_19 sp66_19 sp67_19 11.551961
Rsn66_19 sn66_19 sn67_19 11.551961
Rsp66_20 sp66_20 sp67_20 11.551961
Rsn66_20 sn66_20 sn67_20 11.551961
Rsp66_21 sp66_21 sp67_21 11.551961
Rsn66_21 sn66_21 sn67_21 11.551961
Rsp66_22 sp66_22 sp67_22 11.551961
Rsn66_22 sn66_22 sn67_22 11.551961
Rsp66_23 sp66_23 sp67_23 11.551961
Rsn66_23 sn66_23 sn67_23 11.551961
Rsp66_24 sp66_24 sp67_24 11.551961
Rsn66_24 sn66_24 sn67_24 11.551961
Rsp66_25 sp66_25 sp67_25 11.551961
Rsn66_25 sn66_25 sn67_25 11.551961
Rsp66_26 sp66_26 sp67_26 11.551961
Rsn66_26 sn66_26 sn67_26 11.551961
Rsp66_27 sp66_27 sp67_27 11.551961
Rsn66_27 sn66_27 sn67_27 11.551961
Rsp66_28 sp66_28 sp67_28 11.551961
Rsn66_28 sn66_28 sn67_28 11.551961
Rsp66_29 sp66_29 sp67_29 11.551961
Rsn66_29 sn66_29 sn67_29 11.551961
Rsp66_30 sp66_30 sp67_30 11.551961
Rsn66_30 sn66_30 sn67_30 11.551961
Rsp66_31 sp66_31 sp67_31 11.551961
Rsn66_31 sn66_31 sn67_31 11.551961
Rsp66_32 sp66_32 sp67_32 11.551961
Rsn66_32 sn66_32 sn67_32 11.551961
Rsp66_33 sp66_33 sp67_33 11.551961
Rsn66_33 sn66_33 sn67_33 11.551961
Rsp66_34 sp66_34 sp67_34 11.551961
Rsn66_34 sn66_34 sn67_34 11.551961
Rsp66_35 sp66_35 sp67_35 11.551961
Rsn66_35 sn66_35 sn67_35 11.551961
Rsp66_36 sp66_36 sp67_36 11.551961
Rsn66_36 sn66_36 sn67_36 11.551961
Rsp66_37 sp66_37 sp67_37 11.551961
Rsn66_37 sn66_37 sn67_37 11.551961
Rsp66_38 sp66_38 sp67_38 11.551961
Rsn66_38 sn66_38 sn67_38 11.551961
Rsp66_39 sp66_39 sp67_39 11.551961
Rsn66_39 sn66_39 sn67_39 11.551961
Rsp66_40 sp66_40 sp67_40 11.551961
Rsn66_40 sn66_40 sn67_40 11.551961
Rsp66_41 sp66_41 sp67_41 11.551961
Rsn66_41 sn66_41 sn67_41 11.551961
Rsp66_42 sp66_42 sp67_42 11.551961
Rsn66_42 sn66_42 sn67_42 11.551961
Rsp66_43 sp66_43 sp67_43 11.551961
Rsn66_43 sn66_43 sn67_43 11.551961
Rsp66_44 sp66_44 sp67_44 11.551961
Rsn66_44 sn66_44 sn67_44 11.551961
Rsp66_45 sp66_45 sp67_45 11.551961
Rsn66_45 sn66_45 sn67_45 11.551961
Rsp66_46 sp66_46 sp67_46 11.551961
Rsn66_46 sn66_46 sn67_46 11.551961
Rsp66_47 sp66_47 sp67_47 11.551961
Rsn66_47 sn66_47 sn67_47 11.551961
Rsp66_48 sp66_48 sp67_48 11.551961
Rsn66_48 sn66_48 sn67_48 11.551961
Rsp66_49 sp66_49 sp67_49 11.551961
Rsn66_49 sn66_49 sn67_49 11.551961
Rsp66_50 sp66_50 sp67_50 11.551961
Rsn66_50 sn66_50 sn67_50 11.551961
Rsp66_51 sp66_51 sp67_51 11.551961
Rsn66_51 sn66_51 sn67_51 11.551961
Rsp66_52 sp66_52 sp67_52 11.551961
Rsn66_52 sn66_52 sn67_52 11.551961
Rsp66_53 sp66_53 sp67_53 11.551961
Rsn66_53 sn66_53 sn67_53 11.551961
Rsp66_54 sp66_54 sp67_54 11.551961
Rsn66_54 sn66_54 sn67_54 11.551961
Rsp66_55 sp66_55 sp67_55 11.551961
Rsn66_55 sn66_55 sn67_55 11.551961
Rsp66_56 sp66_56 sp67_56 11.551961
Rsn66_56 sn66_56 sn67_56 11.551961
Rsp66_57 sp66_57 sp67_57 11.551961
Rsn66_57 sn66_57 sn67_57 11.551961
Rsp66_58 sp66_58 sp67_58 11.551961
Rsn66_58 sn66_58 sn67_58 11.551961
Rsp66_59 sp66_59 sp67_59 11.551961
Rsn66_59 sn66_59 sn67_59 11.551961
Rsp66_60 sp66_60 sp67_60 11.551961
Rsn66_60 sn66_60 sn67_60 11.551961
Rsp66_61 sp66_61 sp67_61 11.551961
Rsn66_61 sn66_61 sn67_61 11.551961
Rsp66_62 sp66_62 sp67_62 11.551961
Rsn66_62 sn66_62 sn67_62 11.551961
Rsp66_63 sp66_63 sp67_63 11.551961
Rsn66_63 sn66_63 sn67_63 11.551961
Rsp66_64 sp66_64 sp67_64 11.551961
Rsn66_64 sn66_64 sn67_64 11.551961
Rsp66_65 sp66_65 sp67_65 11.551961
Rsn66_65 sn66_65 sn67_65 11.551961
Rsp66_66 sp66_66 sp67_66 11.551961
Rsn66_66 sn66_66 sn67_66 11.551961
Rsp66_67 sp66_67 sp67_67 11.551961
Rsn66_67 sn66_67 sn67_67 11.551961
Rsp66_68 sp66_68 sp67_68 11.551961
Rsn66_68 sn66_68 sn67_68 11.551961
Rsp66_69 sp66_69 sp67_69 11.551961
Rsn66_69 sn66_69 sn67_69 11.551961
Rsp66_70 sp66_70 sp67_70 11.551961
Rsn66_70 sn66_70 sn67_70 11.551961
Rsp66_71 sp66_71 sp67_71 11.551961
Rsn66_71 sn66_71 sn67_71 11.551961
Rsp66_72 sp66_72 sp67_72 11.551961
Rsn66_72 sn66_72 sn67_72 11.551961
Rsp66_73 sp66_73 sp67_73 11.551961
Rsn66_73 sn66_73 sn67_73 11.551961
Rsp66_74 sp66_74 sp67_74 11.551961
Rsn66_74 sn66_74 sn67_74 11.551961
Rsp66_75 sp66_75 sp67_75 11.551961
Rsn66_75 sn66_75 sn67_75 11.551961
Rsp66_76 sp66_76 sp67_76 11.551961
Rsn66_76 sn66_76 sn67_76 11.551961
Rsp66_77 sp66_77 sp67_77 11.551961
Rsn66_77 sn66_77 sn67_77 11.551961
Rsp66_78 sp66_78 sp67_78 11.551961
Rsn66_78 sn66_78 sn67_78 11.551961
Rsp66_79 sp66_79 sp67_79 11.551961
Rsn66_79 sn66_79 sn67_79 11.551961
Rsp66_80 sp66_80 sp67_80 11.551961
Rsn66_80 sn66_80 sn67_80 11.551961
Rsp66_81 sp66_81 sp67_81 11.551961
Rsn66_81 sn66_81 sn67_81 11.551961
Rsp66_82 sp66_82 sp67_82 11.551961
Rsn66_82 sn66_82 sn67_82 11.551961
Rsp66_83 sp66_83 sp67_83 11.551961
Rsn66_83 sn66_83 sn67_83 11.551961
Rsp66_84 sp66_84 sp67_84 11.551961
Rsn66_84 sn66_84 sn67_84 11.551961
Rsp67_1 sp67_1 sp68_1 11.551961
Rsn67_1 sn67_1 sn68_1 11.551961
Rsp67_2 sp67_2 sp68_2 11.551961
Rsn67_2 sn67_2 sn68_2 11.551961
Rsp67_3 sp67_3 sp68_3 11.551961
Rsn67_3 sn67_3 sn68_3 11.551961
Rsp67_4 sp67_4 sp68_4 11.551961
Rsn67_4 sn67_4 sn68_4 11.551961
Rsp67_5 sp67_5 sp68_5 11.551961
Rsn67_5 sn67_5 sn68_5 11.551961
Rsp67_6 sp67_6 sp68_6 11.551961
Rsn67_6 sn67_6 sn68_6 11.551961
Rsp67_7 sp67_7 sp68_7 11.551961
Rsn67_7 sn67_7 sn68_7 11.551961
Rsp67_8 sp67_8 sp68_8 11.551961
Rsn67_8 sn67_8 sn68_8 11.551961
Rsp67_9 sp67_9 sp68_9 11.551961
Rsn67_9 sn67_9 sn68_9 11.551961
Rsp67_10 sp67_10 sp68_10 11.551961
Rsn67_10 sn67_10 sn68_10 11.551961
Rsp67_11 sp67_11 sp68_11 11.551961
Rsn67_11 sn67_11 sn68_11 11.551961
Rsp67_12 sp67_12 sp68_12 11.551961
Rsn67_12 sn67_12 sn68_12 11.551961
Rsp67_13 sp67_13 sp68_13 11.551961
Rsn67_13 sn67_13 sn68_13 11.551961
Rsp67_14 sp67_14 sp68_14 11.551961
Rsn67_14 sn67_14 sn68_14 11.551961
Rsp67_15 sp67_15 sp68_15 11.551961
Rsn67_15 sn67_15 sn68_15 11.551961
Rsp67_16 sp67_16 sp68_16 11.551961
Rsn67_16 sn67_16 sn68_16 11.551961
Rsp67_17 sp67_17 sp68_17 11.551961
Rsn67_17 sn67_17 sn68_17 11.551961
Rsp67_18 sp67_18 sp68_18 11.551961
Rsn67_18 sn67_18 sn68_18 11.551961
Rsp67_19 sp67_19 sp68_19 11.551961
Rsn67_19 sn67_19 sn68_19 11.551961
Rsp67_20 sp67_20 sp68_20 11.551961
Rsn67_20 sn67_20 sn68_20 11.551961
Rsp67_21 sp67_21 sp68_21 11.551961
Rsn67_21 sn67_21 sn68_21 11.551961
Rsp67_22 sp67_22 sp68_22 11.551961
Rsn67_22 sn67_22 sn68_22 11.551961
Rsp67_23 sp67_23 sp68_23 11.551961
Rsn67_23 sn67_23 sn68_23 11.551961
Rsp67_24 sp67_24 sp68_24 11.551961
Rsn67_24 sn67_24 sn68_24 11.551961
Rsp67_25 sp67_25 sp68_25 11.551961
Rsn67_25 sn67_25 sn68_25 11.551961
Rsp67_26 sp67_26 sp68_26 11.551961
Rsn67_26 sn67_26 sn68_26 11.551961
Rsp67_27 sp67_27 sp68_27 11.551961
Rsn67_27 sn67_27 sn68_27 11.551961
Rsp67_28 sp67_28 sp68_28 11.551961
Rsn67_28 sn67_28 sn68_28 11.551961
Rsp67_29 sp67_29 sp68_29 11.551961
Rsn67_29 sn67_29 sn68_29 11.551961
Rsp67_30 sp67_30 sp68_30 11.551961
Rsn67_30 sn67_30 sn68_30 11.551961
Rsp67_31 sp67_31 sp68_31 11.551961
Rsn67_31 sn67_31 sn68_31 11.551961
Rsp67_32 sp67_32 sp68_32 11.551961
Rsn67_32 sn67_32 sn68_32 11.551961
Rsp67_33 sp67_33 sp68_33 11.551961
Rsn67_33 sn67_33 sn68_33 11.551961
Rsp67_34 sp67_34 sp68_34 11.551961
Rsn67_34 sn67_34 sn68_34 11.551961
Rsp67_35 sp67_35 sp68_35 11.551961
Rsn67_35 sn67_35 sn68_35 11.551961
Rsp67_36 sp67_36 sp68_36 11.551961
Rsn67_36 sn67_36 sn68_36 11.551961
Rsp67_37 sp67_37 sp68_37 11.551961
Rsn67_37 sn67_37 sn68_37 11.551961
Rsp67_38 sp67_38 sp68_38 11.551961
Rsn67_38 sn67_38 sn68_38 11.551961
Rsp67_39 sp67_39 sp68_39 11.551961
Rsn67_39 sn67_39 sn68_39 11.551961
Rsp67_40 sp67_40 sp68_40 11.551961
Rsn67_40 sn67_40 sn68_40 11.551961
Rsp67_41 sp67_41 sp68_41 11.551961
Rsn67_41 sn67_41 sn68_41 11.551961
Rsp67_42 sp67_42 sp68_42 11.551961
Rsn67_42 sn67_42 sn68_42 11.551961
Rsp67_43 sp67_43 sp68_43 11.551961
Rsn67_43 sn67_43 sn68_43 11.551961
Rsp67_44 sp67_44 sp68_44 11.551961
Rsn67_44 sn67_44 sn68_44 11.551961
Rsp67_45 sp67_45 sp68_45 11.551961
Rsn67_45 sn67_45 sn68_45 11.551961
Rsp67_46 sp67_46 sp68_46 11.551961
Rsn67_46 sn67_46 sn68_46 11.551961
Rsp67_47 sp67_47 sp68_47 11.551961
Rsn67_47 sn67_47 sn68_47 11.551961
Rsp67_48 sp67_48 sp68_48 11.551961
Rsn67_48 sn67_48 sn68_48 11.551961
Rsp67_49 sp67_49 sp68_49 11.551961
Rsn67_49 sn67_49 sn68_49 11.551961
Rsp67_50 sp67_50 sp68_50 11.551961
Rsn67_50 sn67_50 sn68_50 11.551961
Rsp67_51 sp67_51 sp68_51 11.551961
Rsn67_51 sn67_51 sn68_51 11.551961
Rsp67_52 sp67_52 sp68_52 11.551961
Rsn67_52 sn67_52 sn68_52 11.551961
Rsp67_53 sp67_53 sp68_53 11.551961
Rsn67_53 sn67_53 sn68_53 11.551961
Rsp67_54 sp67_54 sp68_54 11.551961
Rsn67_54 sn67_54 sn68_54 11.551961
Rsp67_55 sp67_55 sp68_55 11.551961
Rsn67_55 sn67_55 sn68_55 11.551961
Rsp67_56 sp67_56 sp68_56 11.551961
Rsn67_56 sn67_56 sn68_56 11.551961
Rsp67_57 sp67_57 sp68_57 11.551961
Rsn67_57 sn67_57 sn68_57 11.551961
Rsp67_58 sp67_58 sp68_58 11.551961
Rsn67_58 sn67_58 sn68_58 11.551961
Rsp67_59 sp67_59 sp68_59 11.551961
Rsn67_59 sn67_59 sn68_59 11.551961
Rsp67_60 sp67_60 sp68_60 11.551961
Rsn67_60 sn67_60 sn68_60 11.551961
Rsp67_61 sp67_61 sp68_61 11.551961
Rsn67_61 sn67_61 sn68_61 11.551961
Rsp67_62 sp67_62 sp68_62 11.551961
Rsn67_62 sn67_62 sn68_62 11.551961
Rsp67_63 sp67_63 sp68_63 11.551961
Rsn67_63 sn67_63 sn68_63 11.551961
Rsp67_64 sp67_64 sp68_64 11.551961
Rsn67_64 sn67_64 sn68_64 11.551961
Rsp67_65 sp67_65 sp68_65 11.551961
Rsn67_65 sn67_65 sn68_65 11.551961
Rsp67_66 sp67_66 sp68_66 11.551961
Rsn67_66 sn67_66 sn68_66 11.551961
Rsp67_67 sp67_67 sp68_67 11.551961
Rsn67_67 sn67_67 sn68_67 11.551961
Rsp67_68 sp67_68 sp68_68 11.551961
Rsn67_68 sn67_68 sn68_68 11.551961
Rsp67_69 sp67_69 sp68_69 11.551961
Rsn67_69 sn67_69 sn68_69 11.551961
Rsp67_70 sp67_70 sp68_70 11.551961
Rsn67_70 sn67_70 sn68_70 11.551961
Rsp67_71 sp67_71 sp68_71 11.551961
Rsn67_71 sn67_71 sn68_71 11.551961
Rsp67_72 sp67_72 sp68_72 11.551961
Rsn67_72 sn67_72 sn68_72 11.551961
Rsp67_73 sp67_73 sp68_73 11.551961
Rsn67_73 sn67_73 sn68_73 11.551961
Rsp67_74 sp67_74 sp68_74 11.551961
Rsn67_74 sn67_74 sn68_74 11.551961
Rsp67_75 sp67_75 sp68_75 11.551961
Rsn67_75 sn67_75 sn68_75 11.551961
Rsp67_76 sp67_76 sp68_76 11.551961
Rsn67_76 sn67_76 sn68_76 11.551961
Rsp67_77 sp67_77 sp68_77 11.551961
Rsn67_77 sn67_77 sn68_77 11.551961
Rsp67_78 sp67_78 sp68_78 11.551961
Rsn67_78 sn67_78 sn68_78 11.551961
Rsp67_79 sp67_79 sp68_79 11.551961
Rsn67_79 sn67_79 sn68_79 11.551961
Rsp67_80 sp67_80 sp68_80 11.551961
Rsn67_80 sn67_80 sn68_80 11.551961
Rsp67_81 sp67_81 sp68_81 11.551961
Rsn67_81 sn67_81 sn68_81 11.551961
Rsp67_82 sp67_82 sp68_82 11.551961
Rsn67_82 sn67_82 sn68_82 11.551961
Rsp67_83 sp67_83 sp68_83 11.551961
Rsn67_83 sn67_83 sn68_83 11.551961
Rsp67_84 sp67_84 sp68_84 11.551961
Rsn67_84 sn67_84 sn68_84 11.551961
Rsp68_1 sp68_1 sp69_1 11.551961
Rsn68_1 sn68_1 sn69_1 11.551961
Rsp68_2 sp68_2 sp69_2 11.551961
Rsn68_2 sn68_2 sn69_2 11.551961
Rsp68_3 sp68_3 sp69_3 11.551961
Rsn68_3 sn68_3 sn69_3 11.551961
Rsp68_4 sp68_4 sp69_4 11.551961
Rsn68_4 sn68_4 sn69_4 11.551961
Rsp68_5 sp68_5 sp69_5 11.551961
Rsn68_5 sn68_5 sn69_5 11.551961
Rsp68_6 sp68_6 sp69_6 11.551961
Rsn68_6 sn68_6 sn69_6 11.551961
Rsp68_7 sp68_7 sp69_7 11.551961
Rsn68_7 sn68_7 sn69_7 11.551961
Rsp68_8 sp68_8 sp69_8 11.551961
Rsn68_8 sn68_8 sn69_8 11.551961
Rsp68_9 sp68_9 sp69_9 11.551961
Rsn68_9 sn68_9 sn69_9 11.551961
Rsp68_10 sp68_10 sp69_10 11.551961
Rsn68_10 sn68_10 sn69_10 11.551961
Rsp68_11 sp68_11 sp69_11 11.551961
Rsn68_11 sn68_11 sn69_11 11.551961
Rsp68_12 sp68_12 sp69_12 11.551961
Rsn68_12 sn68_12 sn69_12 11.551961
Rsp68_13 sp68_13 sp69_13 11.551961
Rsn68_13 sn68_13 sn69_13 11.551961
Rsp68_14 sp68_14 sp69_14 11.551961
Rsn68_14 sn68_14 sn69_14 11.551961
Rsp68_15 sp68_15 sp69_15 11.551961
Rsn68_15 sn68_15 sn69_15 11.551961
Rsp68_16 sp68_16 sp69_16 11.551961
Rsn68_16 sn68_16 sn69_16 11.551961
Rsp68_17 sp68_17 sp69_17 11.551961
Rsn68_17 sn68_17 sn69_17 11.551961
Rsp68_18 sp68_18 sp69_18 11.551961
Rsn68_18 sn68_18 sn69_18 11.551961
Rsp68_19 sp68_19 sp69_19 11.551961
Rsn68_19 sn68_19 sn69_19 11.551961
Rsp68_20 sp68_20 sp69_20 11.551961
Rsn68_20 sn68_20 sn69_20 11.551961
Rsp68_21 sp68_21 sp69_21 11.551961
Rsn68_21 sn68_21 sn69_21 11.551961
Rsp68_22 sp68_22 sp69_22 11.551961
Rsn68_22 sn68_22 sn69_22 11.551961
Rsp68_23 sp68_23 sp69_23 11.551961
Rsn68_23 sn68_23 sn69_23 11.551961
Rsp68_24 sp68_24 sp69_24 11.551961
Rsn68_24 sn68_24 sn69_24 11.551961
Rsp68_25 sp68_25 sp69_25 11.551961
Rsn68_25 sn68_25 sn69_25 11.551961
Rsp68_26 sp68_26 sp69_26 11.551961
Rsn68_26 sn68_26 sn69_26 11.551961
Rsp68_27 sp68_27 sp69_27 11.551961
Rsn68_27 sn68_27 sn69_27 11.551961
Rsp68_28 sp68_28 sp69_28 11.551961
Rsn68_28 sn68_28 sn69_28 11.551961
Rsp68_29 sp68_29 sp69_29 11.551961
Rsn68_29 sn68_29 sn69_29 11.551961
Rsp68_30 sp68_30 sp69_30 11.551961
Rsn68_30 sn68_30 sn69_30 11.551961
Rsp68_31 sp68_31 sp69_31 11.551961
Rsn68_31 sn68_31 sn69_31 11.551961
Rsp68_32 sp68_32 sp69_32 11.551961
Rsn68_32 sn68_32 sn69_32 11.551961
Rsp68_33 sp68_33 sp69_33 11.551961
Rsn68_33 sn68_33 sn69_33 11.551961
Rsp68_34 sp68_34 sp69_34 11.551961
Rsn68_34 sn68_34 sn69_34 11.551961
Rsp68_35 sp68_35 sp69_35 11.551961
Rsn68_35 sn68_35 sn69_35 11.551961
Rsp68_36 sp68_36 sp69_36 11.551961
Rsn68_36 sn68_36 sn69_36 11.551961
Rsp68_37 sp68_37 sp69_37 11.551961
Rsn68_37 sn68_37 sn69_37 11.551961
Rsp68_38 sp68_38 sp69_38 11.551961
Rsn68_38 sn68_38 sn69_38 11.551961
Rsp68_39 sp68_39 sp69_39 11.551961
Rsn68_39 sn68_39 sn69_39 11.551961
Rsp68_40 sp68_40 sp69_40 11.551961
Rsn68_40 sn68_40 sn69_40 11.551961
Rsp68_41 sp68_41 sp69_41 11.551961
Rsn68_41 sn68_41 sn69_41 11.551961
Rsp68_42 sp68_42 sp69_42 11.551961
Rsn68_42 sn68_42 sn69_42 11.551961
Rsp68_43 sp68_43 sp69_43 11.551961
Rsn68_43 sn68_43 sn69_43 11.551961
Rsp68_44 sp68_44 sp69_44 11.551961
Rsn68_44 sn68_44 sn69_44 11.551961
Rsp68_45 sp68_45 sp69_45 11.551961
Rsn68_45 sn68_45 sn69_45 11.551961
Rsp68_46 sp68_46 sp69_46 11.551961
Rsn68_46 sn68_46 sn69_46 11.551961
Rsp68_47 sp68_47 sp69_47 11.551961
Rsn68_47 sn68_47 sn69_47 11.551961
Rsp68_48 sp68_48 sp69_48 11.551961
Rsn68_48 sn68_48 sn69_48 11.551961
Rsp68_49 sp68_49 sp69_49 11.551961
Rsn68_49 sn68_49 sn69_49 11.551961
Rsp68_50 sp68_50 sp69_50 11.551961
Rsn68_50 sn68_50 sn69_50 11.551961
Rsp68_51 sp68_51 sp69_51 11.551961
Rsn68_51 sn68_51 sn69_51 11.551961
Rsp68_52 sp68_52 sp69_52 11.551961
Rsn68_52 sn68_52 sn69_52 11.551961
Rsp68_53 sp68_53 sp69_53 11.551961
Rsn68_53 sn68_53 sn69_53 11.551961
Rsp68_54 sp68_54 sp69_54 11.551961
Rsn68_54 sn68_54 sn69_54 11.551961
Rsp68_55 sp68_55 sp69_55 11.551961
Rsn68_55 sn68_55 sn69_55 11.551961
Rsp68_56 sp68_56 sp69_56 11.551961
Rsn68_56 sn68_56 sn69_56 11.551961
Rsp68_57 sp68_57 sp69_57 11.551961
Rsn68_57 sn68_57 sn69_57 11.551961
Rsp68_58 sp68_58 sp69_58 11.551961
Rsn68_58 sn68_58 sn69_58 11.551961
Rsp68_59 sp68_59 sp69_59 11.551961
Rsn68_59 sn68_59 sn69_59 11.551961
Rsp68_60 sp68_60 sp69_60 11.551961
Rsn68_60 sn68_60 sn69_60 11.551961
Rsp68_61 sp68_61 sp69_61 11.551961
Rsn68_61 sn68_61 sn69_61 11.551961
Rsp68_62 sp68_62 sp69_62 11.551961
Rsn68_62 sn68_62 sn69_62 11.551961
Rsp68_63 sp68_63 sp69_63 11.551961
Rsn68_63 sn68_63 sn69_63 11.551961
Rsp68_64 sp68_64 sp69_64 11.551961
Rsn68_64 sn68_64 sn69_64 11.551961
Rsp68_65 sp68_65 sp69_65 11.551961
Rsn68_65 sn68_65 sn69_65 11.551961
Rsp68_66 sp68_66 sp69_66 11.551961
Rsn68_66 sn68_66 sn69_66 11.551961
Rsp68_67 sp68_67 sp69_67 11.551961
Rsn68_67 sn68_67 sn69_67 11.551961
Rsp68_68 sp68_68 sp69_68 11.551961
Rsn68_68 sn68_68 sn69_68 11.551961
Rsp68_69 sp68_69 sp69_69 11.551961
Rsn68_69 sn68_69 sn69_69 11.551961
Rsp68_70 sp68_70 sp69_70 11.551961
Rsn68_70 sn68_70 sn69_70 11.551961
Rsp68_71 sp68_71 sp69_71 11.551961
Rsn68_71 sn68_71 sn69_71 11.551961
Rsp68_72 sp68_72 sp69_72 11.551961
Rsn68_72 sn68_72 sn69_72 11.551961
Rsp68_73 sp68_73 sp69_73 11.551961
Rsn68_73 sn68_73 sn69_73 11.551961
Rsp68_74 sp68_74 sp69_74 11.551961
Rsn68_74 sn68_74 sn69_74 11.551961
Rsp68_75 sp68_75 sp69_75 11.551961
Rsn68_75 sn68_75 sn69_75 11.551961
Rsp68_76 sp68_76 sp69_76 11.551961
Rsn68_76 sn68_76 sn69_76 11.551961
Rsp68_77 sp68_77 sp69_77 11.551961
Rsn68_77 sn68_77 sn69_77 11.551961
Rsp68_78 sp68_78 sp69_78 11.551961
Rsn68_78 sn68_78 sn69_78 11.551961
Rsp68_79 sp68_79 sp69_79 11.551961
Rsn68_79 sn68_79 sn69_79 11.551961
Rsp68_80 sp68_80 sp69_80 11.551961
Rsn68_80 sn68_80 sn69_80 11.551961
Rsp68_81 sp68_81 sp69_81 11.551961
Rsn68_81 sn68_81 sn69_81 11.551961
Rsp68_82 sp68_82 sp69_82 11.551961
Rsn68_82 sn68_82 sn69_82 11.551961
Rsp68_83 sp68_83 sp69_83 11.551961
Rsn68_83 sn68_83 sn69_83 11.551961
Rsp68_84 sp68_84 sp69_84 11.551961
Rsn68_84 sn68_84 sn69_84 11.551961
Rsp69_1 sp69_1 sp70_1 11.551961
Rsn69_1 sn69_1 sn70_1 11.551961
Rsp69_2 sp69_2 sp70_2 11.551961
Rsn69_2 sn69_2 sn70_2 11.551961
Rsp69_3 sp69_3 sp70_3 11.551961
Rsn69_3 sn69_3 sn70_3 11.551961
Rsp69_4 sp69_4 sp70_4 11.551961
Rsn69_4 sn69_4 sn70_4 11.551961
Rsp69_5 sp69_5 sp70_5 11.551961
Rsn69_5 sn69_5 sn70_5 11.551961
Rsp69_6 sp69_6 sp70_6 11.551961
Rsn69_6 sn69_6 sn70_6 11.551961
Rsp69_7 sp69_7 sp70_7 11.551961
Rsn69_7 sn69_7 sn70_7 11.551961
Rsp69_8 sp69_8 sp70_8 11.551961
Rsn69_8 sn69_8 sn70_8 11.551961
Rsp69_9 sp69_9 sp70_9 11.551961
Rsn69_9 sn69_9 sn70_9 11.551961
Rsp69_10 sp69_10 sp70_10 11.551961
Rsn69_10 sn69_10 sn70_10 11.551961
Rsp69_11 sp69_11 sp70_11 11.551961
Rsn69_11 sn69_11 sn70_11 11.551961
Rsp69_12 sp69_12 sp70_12 11.551961
Rsn69_12 sn69_12 sn70_12 11.551961
Rsp69_13 sp69_13 sp70_13 11.551961
Rsn69_13 sn69_13 sn70_13 11.551961
Rsp69_14 sp69_14 sp70_14 11.551961
Rsn69_14 sn69_14 sn70_14 11.551961
Rsp69_15 sp69_15 sp70_15 11.551961
Rsn69_15 sn69_15 sn70_15 11.551961
Rsp69_16 sp69_16 sp70_16 11.551961
Rsn69_16 sn69_16 sn70_16 11.551961
Rsp69_17 sp69_17 sp70_17 11.551961
Rsn69_17 sn69_17 sn70_17 11.551961
Rsp69_18 sp69_18 sp70_18 11.551961
Rsn69_18 sn69_18 sn70_18 11.551961
Rsp69_19 sp69_19 sp70_19 11.551961
Rsn69_19 sn69_19 sn70_19 11.551961
Rsp69_20 sp69_20 sp70_20 11.551961
Rsn69_20 sn69_20 sn70_20 11.551961
Rsp69_21 sp69_21 sp70_21 11.551961
Rsn69_21 sn69_21 sn70_21 11.551961
Rsp69_22 sp69_22 sp70_22 11.551961
Rsn69_22 sn69_22 sn70_22 11.551961
Rsp69_23 sp69_23 sp70_23 11.551961
Rsn69_23 sn69_23 sn70_23 11.551961
Rsp69_24 sp69_24 sp70_24 11.551961
Rsn69_24 sn69_24 sn70_24 11.551961
Rsp69_25 sp69_25 sp70_25 11.551961
Rsn69_25 sn69_25 sn70_25 11.551961
Rsp69_26 sp69_26 sp70_26 11.551961
Rsn69_26 sn69_26 sn70_26 11.551961
Rsp69_27 sp69_27 sp70_27 11.551961
Rsn69_27 sn69_27 sn70_27 11.551961
Rsp69_28 sp69_28 sp70_28 11.551961
Rsn69_28 sn69_28 sn70_28 11.551961
Rsp69_29 sp69_29 sp70_29 11.551961
Rsn69_29 sn69_29 sn70_29 11.551961
Rsp69_30 sp69_30 sp70_30 11.551961
Rsn69_30 sn69_30 sn70_30 11.551961
Rsp69_31 sp69_31 sp70_31 11.551961
Rsn69_31 sn69_31 sn70_31 11.551961
Rsp69_32 sp69_32 sp70_32 11.551961
Rsn69_32 sn69_32 sn70_32 11.551961
Rsp69_33 sp69_33 sp70_33 11.551961
Rsn69_33 sn69_33 sn70_33 11.551961
Rsp69_34 sp69_34 sp70_34 11.551961
Rsn69_34 sn69_34 sn70_34 11.551961
Rsp69_35 sp69_35 sp70_35 11.551961
Rsn69_35 sn69_35 sn70_35 11.551961
Rsp69_36 sp69_36 sp70_36 11.551961
Rsn69_36 sn69_36 sn70_36 11.551961
Rsp69_37 sp69_37 sp70_37 11.551961
Rsn69_37 sn69_37 sn70_37 11.551961
Rsp69_38 sp69_38 sp70_38 11.551961
Rsn69_38 sn69_38 sn70_38 11.551961
Rsp69_39 sp69_39 sp70_39 11.551961
Rsn69_39 sn69_39 sn70_39 11.551961
Rsp69_40 sp69_40 sp70_40 11.551961
Rsn69_40 sn69_40 sn70_40 11.551961
Rsp69_41 sp69_41 sp70_41 11.551961
Rsn69_41 sn69_41 sn70_41 11.551961
Rsp69_42 sp69_42 sp70_42 11.551961
Rsn69_42 sn69_42 sn70_42 11.551961
Rsp69_43 sp69_43 sp70_43 11.551961
Rsn69_43 sn69_43 sn70_43 11.551961
Rsp69_44 sp69_44 sp70_44 11.551961
Rsn69_44 sn69_44 sn70_44 11.551961
Rsp69_45 sp69_45 sp70_45 11.551961
Rsn69_45 sn69_45 sn70_45 11.551961
Rsp69_46 sp69_46 sp70_46 11.551961
Rsn69_46 sn69_46 sn70_46 11.551961
Rsp69_47 sp69_47 sp70_47 11.551961
Rsn69_47 sn69_47 sn70_47 11.551961
Rsp69_48 sp69_48 sp70_48 11.551961
Rsn69_48 sn69_48 sn70_48 11.551961
Rsp69_49 sp69_49 sp70_49 11.551961
Rsn69_49 sn69_49 sn70_49 11.551961
Rsp69_50 sp69_50 sp70_50 11.551961
Rsn69_50 sn69_50 sn70_50 11.551961
Rsp69_51 sp69_51 sp70_51 11.551961
Rsn69_51 sn69_51 sn70_51 11.551961
Rsp69_52 sp69_52 sp70_52 11.551961
Rsn69_52 sn69_52 sn70_52 11.551961
Rsp69_53 sp69_53 sp70_53 11.551961
Rsn69_53 sn69_53 sn70_53 11.551961
Rsp69_54 sp69_54 sp70_54 11.551961
Rsn69_54 sn69_54 sn70_54 11.551961
Rsp69_55 sp69_55 sp70_55 11.551961
Rsn69_55 sn69_55 sn70_55 11.551961
Rsp69_56 sp69_56 sp70_56 11.551961
Rsn69_56 sn69_56 sn70_56 11.551961
Rsp69_57 sp69_57 sp70_57 11.551961
Rsn69_57 sn69_57 sn70_57 11.551961
Rsp69_58 sp69_58 sp70_58 11.551961
Rsn69_58 sn69_58 sn70_58 11.551961
Rsp69_59 sp69_59 sp70_59 11.551961
Rsn69_59 sn69_59 sn70_59 11.551961
Rsp69_60 sp69_60 sp70_60 11.551961
Rsn69_60 sn69_60 sn70_60 11.551961
Rsp69_61 sp69_61 sp70_61 11.551961
Rsn69_61 sn69_61 sn70_61 11.551961
Rsp69_62 sp69_62 sp70_62 11.551961
Rsn69_62 sn69_62 sn70_62 11.551961
Rsp69_63 sp69_63 sp70_63 11.551961
Rsn69_63 sn69_63 sn70_63 11.551961
Rsp69_64 sp69_64 sp70_64 11.551961
Rsn69_64 sn69_64 sn70_64 11.551961
Rsp69_65 sp69_65 sp70_65 11.551961
Rsn69_65 sn69_65 sn70_65 11.551961
Rsp69_66 sp69_66 sp70_66 11.551961
Rsn69_66 sn69_66 sn70_66 11.551961
Rsp69_67 sp69_67 sp70_67 11.551961
Rsn69_67 sn69_67 sn70_67 11.551961
Rsp69_68 sp69_68 sp70_68 11.551961
Rsn69_68 sn69_68 sn70_68 11.551961
Rsp69_69 sp69_69 sp70_69 11.551961
Rsn69_69 sn69_69 sn70_69 11.551961
Rsp69_70 sp69_70 sp70_70 11.551961
Rsn69_70 sn69_70 sn70_70 11.551961
Rsp69_71 sp69_71 sp70_71 11.551961
Rsn69_71 sn69_71 sn70_71 11.551961
Rsp69_72 sp69_72 sp70_72 11.551961
Rsn69_72 sn69_72 sn70_72 11.551961
Rsp69_73 sp69_73 sp70_73 11.551961
Rsn69_73 sn69_73 sn70_73 11.551961
Rsp69_74 sp69_74 sp70_74 11.551961
Rsn69_74 sn69_74 sn70_74 11.551961
Rsp69_75 sp69_75 sp70_75 11.551961
Rsn69_75 sn69_75 sn70_75 11.551961
Rsp69_76 sp69_76 sp70_76 11.551961
Rsn69_76 sn69_76 sn70_76 11.551961
Rsp69_77 sp69_77 sp70_77 11.551961
Rsn69_77 sn69_77 sn70_77 11.551961
Rsp69_78 sp69_78 sp70_78 11.551961
Rsn69_78 sn69_78 sn70_78 11.551961
Rsp69_79 sp69_79 sp70_79 11.551961
Rsn69_79 sn69_79 sn70_79 11.551961
Rsp69_80 sp69_80 sp70_80 11.551961
Rsn69_80 sn69_80 sn70_80 11.551961
Rsp69_81 sp69_81 sp70_81 11.551961
Rsn69_81 sn69_81 sn70_81 11.551961
Rsp69_82 sp69_82 sp70_82 11.551961
Rsn69_82 sn69_82 sn70_82 11.551961
Rsp69_83 sp69_83 sp70_83 11.551961
Rsn69_83 sn69_83 sn70_83 11.551961
Rsp69_84 sp69_84 sp70_84 11.551961
Rsn69_84 sn69_84 sn70_84 11.551961
Rsp70_1 sp70_1 sp71_1 11.551961
Rsn70_1 sn70_1 sn71_1 11.551961
Rsp70_2 sp70_2 sp71_2 11.551961
Rsn70_2 sn70_2 sn71_2 11.551961
Rsp70_3 sp70_3 sp71_3 11.551961
Rsn70_3 sn70_3 sn71_3 11.551961
Rsp70_4 sp70_4 sp71_4 11.551961
Rsn70_4 sn70_4 sn71_4 11.551961
Rsp70_5 sp70_5 sp71_5 11.551961
Rsn70_5 sn70_5 sn71_5 11.551961
Rsp70_6 sp70_6 sp71_6 11.551961
Rsn70_6 sn70_6 sn71_6 11.551961
Rsp70_7 sp70_7 sp71_7 11.551961
Rsn70_7 sn70_7 sn71_7 11.551961
Rsp70_8 sp70_8 sp71_8 11.551961
Rsn70_8 sn70_8 sn71_8 11.551961
Rsp70_9 sp70_9 sp71_9 11.551961
Rsn70_9 sn70_9 sn71_9 11.551961
Rsp70_10 sp70_10 sp71_10 11.551961
Rsn70_10 sn70_10 sn71_10 11.551961
Rsp70_11 sp70_11 sp71_11 11.551961
Rsn70_11 sn70_11 sn71_11 11.551961
Rsp70_12 sp70_12 sp71_12 11.551961
Rsn70_12 sn70_12 sn71_12 11.551961
Rsp70_13 sp70_13 sp71_13 11.551961
Rsn70_13 sn70_13 sn71_13 11.551961
Rsp70_14 sp70_14 sp71_14 11.551961
Rsn70_14 sn70_14 sn71_14 11.551961
Rsp70_15 sp70_15 sp71_15 11.551961
Rsn70_15 sn70_15 sn71_15 11.551961
Rsp70_16 sp70_16 sp71_16 11.551961
Rsn70_16 sn70_16 sn71_16 11.551961
Rsp70_17 sp70_17 sp71_17 11.551961
Rsn70_17 sn70_17 sn71_17 11.551961
Rsp70_18 sp70_18 sp71_18 11.551961
Rsn70_18 sn70_18 sn71_18 11.551961
Rsp70_19 sp70_19 sp71_19 11.551961
Rsn70_19 sn70_19 sn71_19 11.551961
Rsp70_20 sp70_20 sp71_20 11.551961
Rsn70_20 sn70_20 sn71_20 11.551961
Rsp70_21 sp70_21 sp71_21 11.551961
Rsn70_21 sn70_21 sn71_21 11.551961
Rsp70_22 sp70_22 sp71_22 11.551961
Rsn70_22 sn70_22 sn71_22 11.551961
Rsp70_23 sp70_23 sp71_23 11.551961
Rsn70_23 sn70_23 sn71_23 11.551961
Rsp70_24 sp70_24 sp71_24 11.551961
Rsn70_24 sn70_24 sn71_24 11.551961
Rsp70_25 sp70_25 sp71_25 11.551961
Rsn70_25 sn70_25 sn71_25 11.551961
Rsp70_26 sp70_26 sp71_26 11.551961
Rsn70_26 sn70_26 sn71_26 11.551961
Rsp70_27 sp70_27 sp71_27 11.551961
Rsn70_27 sn70_27 sn71_27 11.551961
Rsp70_28 sp70_28 sp71_28 11.551961
Rsn70_28 sn70_28 sn71_28 11.551961
Rsp70_29 sp70_29 sp71_29 11.551961
Rsn70_29 sn70_29 sn71_29 11.551961
Rsp70_30 sp70_30 sp71_30 11.551961
Rsn70_30 sn70_30 sn71_30 11.551961
Rsp70_31 sp70_31 sp71_31 11.551961
Rsn70_31 sn70_31 sn71_31 11.551961
Rsp70_32 sp70_32 sp71_32 11.551961
Rsn70_32 sn70_32 sn71_32 11.551961
Rsp70_33 sp70_33 sp71_33 11.551961
Rsn70_33 sn70_33 sn71_33 11.551961
Rsp70_34 sp70_34 sp71_34 11.551961
Rsn70_34 sn70_34 sn71_34 11.551961
Rsp70_35 sp70_35 sp71_35 11.551961
Rsn70_35 sn70_35 sn71_35 11.551961
Rsp70_36 sp70_36 sp71_36 11.551961
Rsn70_36 sn70_36 sn71_36 11.551961
Rsp70_37 sp70_37 sp71_37 11.551961
Rsn70_37 sn70_37 sn71_37 11.551961
Rsp70_38 sp70_38 sp71_38 11.551961
Rsn70_38 sn70_38 sn71_38 11.551961
Rsp70_39 sp70_39 sp71_39 11.551961
Rsn70_39 sn70_39 sn71_39 11.551961
Rsp70_40 sp70_40 sp71_40 11.551961
Rsn70_40 sn70_40 sn71_40 11.551961
Rsp70_41 sp70_41 sp71_41 11.551961
Rsn70_41 sn70_41 sn71_41 11.551961
Rsp70_42 sp70_42 sp71_42 11.551961
Rsn70_42 sn70_42 sn71_42 11.551961
Rsp70_43 sp70_43 sp71_43 11.551961
Rsn70_43 sn70_43 sn71_43 11.551961
Rsp70_44 sp70_44 sp71_44 11.551961
Rsn70_44 sn70_44 sn71_44 11.551961
Rsp70_45 sp70_45 sp71_45 11.551961
Rsn70_45 sn70_45 sn71_45 11.551961
Rsp70_46 sp70_46 sp71_46 11.551961
Rsn70_46 sn70_46 sn71_46 11.551961
Rsp70_47 sp70_47 sp71_47 11.551961
Rsn70_47 sn70_47 sn71_47 11.551961
Rsp70_48 sp70_48 sp71_48 11.551961
Rsn70_48 sn70_48 sn71_48 11.551961
Rsp70_49 sp70_49 sp71_49 11.551961
Rsn70_49 sn70_49 sn71_49 11.551961
Rsp70_50 sp70_50 sp71_50 11.551961
Rsn70_50 sn70_50 sn71_50 11.551961
Rsp70_51 sp70_51 sp71_51 11.551961
Rsn70_51 sn70_51 sn71_51 11.551961
Rsp70_52 sp70_52 sp71_52 11.551961
Rsn70_52 sn70_52 sn71_52 11.551961
Rsp70_53 sp70_53 sp71_53 11.551961
Rsn70_53 sn70_53 sn71_53 11.551961
Rsp70_54 sp70_54 sp71_54 11.551961
Rsn70_54 sn70_54 sn71_54 11.551961
Rsp70_55 sp70_55 sp71_55 11.551961
Rsn70_55 sn70_55 sn71_55 11.551961
Rsp70_56 sp70_56 sp71_56 11.551961
Rsn70_56 sn70_56 sn71_56 11.551961
Rsp70_57 sp70_57 sp71_57 11.551961
Rsn70_57 sn70_57 sn71_57 11.551961
Rsp70_58 sp70_58 sp71_58 11.551961
Rsn70_58 sn70_58 sn71_58 11.551961
Rsp70_59 sp70_59 sp71_59 11.551961
Rsn70_59 sn70_59 sn71_59 11.551961
Rsp70_60 sp70_60 sp71_60 11.551961
Rsn70_60 sn70_60 sn71_60 11.551961
Rsp70_61 sp70_61 sp71_61 11.551961
Rsn70_61 sn70_61 sn71_61 11.551961
Rsp70_62 sp70_62 sp71_62 11.551961
Rsn70_62 sn70_62 sn71_62 11.551961
Rsp70_63 sp70_63 sp71_63 11.551961
Rsn70_63 sn70_63 sn71_63 11.551961
Rsp70_64 sp70_64 sp71_64 11.551961
Rsn70_64 sn70_64 sn71_64 11.551961
Rsp70_65 sp70_65 sp71_65 11.551961
Rsn70_65 sn70_65 sn71_65 11.551961
Rsp70_66 sp70_66 sp71_66 11.551961
Rsn70_66 sn70_66 sn71_66 11.551961
Rsp70_67 sp70_67 sp71_67 11.551961
Rsn70_67 sn70_67 sn71_67 11.551961
Rsp70_68 sp70_68 sp71_68 11.551961
Rsn70_68 sn70_68 sn71_68 11.551961
Rsp70_69 sp70_69 sp71_69 11.551961
Rsn70_69 sn70_69 sn71_69 11.551961
Rsp70_70 sp70_70 sp71_70 11.551961
Rsn70_70 sn70_70 sn71_70 11.551961
Rsp70_71 sp70_71 sp71_71 11.551961
Rsn70_71 sn70_71 sn71_71 11.551961
Rsp70_72 sp70_72 sp71_72 11.551961
Rsn70_72 sn70_72 sn71_72 11.551961
Rsp70_73 sp70_73 sp71_73 11.551961
Rsn70_73 sn70_73 sn71_73 11.551961
Rsp70_74 sp70_74 sp71_74 11.551961
Rsn70_74 sn70_74 sn71_74 11.551961
Rsp70_75 sp70_75 sp71_75 11.551961
Rsn70_75 sn70_75 sn71_75 11.551961
Rsp70_76 sp70_76 sp71_76 11.551961
Rsn70_76 sn70_76 sn71_76 11.551961
Rsp70_77 sp70_77 sp71_77 11.551961
Rsn70_77 sn70_77 sn71_77 11.551961
Rsp70_78 sp70_78 sp71_78 11.551961
Rsn70_78 sn70_78 sn71_78 11.551961
Rsp70_79 sp70_79 sp71_79 11.551961
Rsn70_79 sn70_79 sn71_79 11.551961
Rsp70_80 sp70_80 sp71_80 11.551961
Rsn70_80 sn70_80 sn71_80 11.551961
Rsp70_81 sp70_81 sp71_81 11.551961
Rsn70_81 sn70_81 sn71_81 11.551961
Rsp70_82 sp70_82 sp71_82 11.551961
Rsn70_82 sn70_82 sn71_82 11.551961
Rsp70_83 sp70_83 sp71_83 11.551961
Rsn70_83 sn70_83 sn71_83 11.551961
Rsp70_84 sp70_84 sp71_84 11.551961
Rsn70_84 sn70_84 sn71_84 11.551961
Rsp71_1 sp71_1 sp72_1 11.551961
Rsn71_1 sn71_1 sn72_1 11.551961
Rsp71_2 sp71_2 sp72_2 11.551961
Rsn71_2 sn71_2 sn72_2 11.551961
Rsp71_3 sp71_3 sp72_3 11.551961
Rsn71_3 sn71_3 sn72_3 11.551961
Rsp71_4 sp71_4 sp72_4 11.551961
Rsn71_4 sn71_4 sn72_4 11.551961
Rsp71_5 sp71_5 sp72_5 11.551961
Rsn71_5 sn71_5 sn72_5 11.551961
Rsp71_6 sp71_6 sp72_6 11.551961
Rsn71_6 sn71_6 sn72_6 11.551961
Rsp71_7 sp71_7 sp72_7 11.551961
Rsn71_7 sn71_7 sn72_7 11.551961
Rsp71_8 sp71_8 sp72_8 11.551961
Rsn71_8 sn71_8 sn72_8 11.551961
Rsp71_9 sp71_9 sp72_9 11.551961
Rsn71_9 sn71_9 sn72_9 11.551961
Rsp71_10 sp71_10 sp72_10 11.551961
Rsn71_10 sn71_10 sn72_10 11.551961
Rsp71_11 sp71_11 sp72_11 11.551961
Rsn71_11 sn71_11 sn72_11 11.551961
Rsp71_12 sp71_12 sp72_12 11.551961
Rsn71_12 sn71_12 sn72_12 11.551961
Rsp71_13 sp71_13 sp72_13 11.551961
Rsn71_13 sn71_13 sn72_13 11.551961
Rsp71_14 sp71_14 sp72_14 11.551961
Rsn71_14 sn71_14 sn72_14 11.551961
Rsp71_15 sp71_15 sp72_15 11.551961
Rsn71_15 sn71_15 sn72_15 11.551961
Rsp71_16 sp71_16 sp72_16 11.551961
Rsn71_16 sn71_16 sn72_16 11.551961
Rsp71_17 sp71_17 sp72_17 11.551961
Rsn71_17 sn71_17 sn72_17 11.551961
Rsp71_18 sp71_18 sp72_18 11.551961
Rsn71_18 sn71_18 sn72_18 11.551961
Rsp71_19 sp71_19 sp72_19 11.551961
Rsn71_19 sn71_19 sn72_19 11.551961
Rsp71_20 sp71_20 sp72_20 11.551961
Rsn71_20 sn71_20 sn72_20 11.551961
Rsp71_21 sp71_21 sp72_21 11.551961
Rsn71_21 sn71_21 sn72_21 11.551961
Rsp71_22 sp71_22 sp72_22 11.551961
Rsn71_22 sn71_22 sn72_22 11.551961
Rsp71_23 sp71_23 sp72_23 11.551961
Rsn71_23 sn71_23 sn72_23 11.551961
Rsp71_24 sp71_24 sp72_24 11.551961
Rsn71_24 sn71_24 sn72_24 11.551961
Rsp71_25 sp71_25 sp72_25 11.551961
Rsn71_25 sn71_25 sn72_25 11.551961
Rsp71_26 sp71_26 sp72_26 11.551961
Rsn71_26 sn71_26 sn72_26 11.551961
Rsp71_27 sp71_27 sp72_27 11.551961
Rsn71_27 sn71_27 sn72_27 11.551961
Rsp71_28 sp71_28 sp72_28 11.551961
Rsn71_28 sn71_28 sn72_28 11.551961
Rsp71_29 sp71_29 sp72_29 11.551961
Rsn71_29 sn71_29 sn72_29 11.551961
Rsp71_30 sp71_30 sp72_30 11.551961
Rsn71_30 sn71_30 sn72_30 11.551961
Rsp71_31 sp71_31 sp72_31 11.551961
Rsn71_31 sn71_31 sn72_31 11.551961
Rsp71_32 sp71_32 sp72_32 11.551961
Rsn71_32 sn71_32 sn72_32 11.551961
Rsp71_33 sp71_33 sp72_33 11.551961
Rsn71_33 sn71_33 sn72_33 11.551961
Rsp71_34 sp71_34 sp72_34 11.551961
Rsn71_34 sn71_34 sn72_34 11.551961
Rsp71_35 sp71_35 sp72_35 11.551961
Rsn71_35 sn71_35 sn72_35 11.551961
Rsp71_36 sp71_36 sp72_36 11.551961
Rsn71_36 sn71_36 sn72_36 11.551961
Rsp71_37 sp71_37 sp72_37 11.551961
Rsn71_37 sn71_37 sn72_37 11.551961
Rsp71_38 sp71_38 sp72_38 11.551961
Rsn71_38 sn71_38 sn72_38 11.551961
Rsp71_39 sp71_39 sp72_39 11.551961
Rsn71_39 sn71_39 sn72_39 11.551961
Rsp71_40 sp71_40 sp72_40 11.551961
Rsn71_40 sn71_40 sn72_40 11.551961
Rsp71_41 sp71_41 sp72_41 11.551961
Rsn71_41 sn71_41 sn72_41 11.551961
Rsp71_42 sp71_42 sp72_42 11.551961
Rsn71_42 sn71_42 sn72_42 11.551961
Rsp71_43 sp71_43 sp72_43 11.551961
Rsn71_43 sn71_43 sn72_43 11.551961
Rsp71_44 sp71_44 sp72_44 11.551961
Rsn71_44 sn71_44 sn72_44 11.551961
Rsp71_45 sp71_45 sp72_45 11.551961
Rsn71_45 sn71_45 sn72_45 11.551961
Rsp71_46 sp71_46 sp72_46 11.551961
Rsn71_46 sn71_46 sn72_46 11.551961
Rsp71_47 sp71_47 sp72_47 11.551961
Rsn71_47 sn71_47 sn72_47 11.551961
Rsp71_48 sp71_48 sp72_48 11.551961
Rsn71_48 sn71_48 sn72_48 11.551961
Rsp71_49 sp71_49 sp72_49 11.551961
Rsn71_49 sn71_49 sn72_49 11.551961
Rsp71_50 sp71_50 sp72_50 11.551961
Rsn71_50 sn71_50 sn72_50 11.551961
Rsp71_51 sp71_51 sp72_51 11.551961
Rsn71_51 sn71_51 sn72_51 11.551961
Rsp71_52 sp71_52 sp72_52 11.551961
Rsn71_52 sn71_52 sn72_52 11.551961
Rsp71_53 sp71_53 sp72_53 11.551961
Rsn71_53 sn71_53 sn72_53 11.551961
Rsp71_54 sp71_54 sp72_54 11.551961
Rsn71_54 sn71_54 sn72_54 11.551961
Rsp71_55 sp71_55 sp72_55 11.551961
Rsn71_55 sn71_55 sn72_55 11.551961
Rsp71_56 sp71_56 sp72_56 11.551961
Rsn71_56 sn71_56 sn72_56 11.551961
Rsp71_57 sp71_57 sp72_57 11.551961
Rsn71_57 sn71_57 sn72_57 11.551961
Rsp71_58 sp71_58 sp72_58 11.551961
Rsn71_58 sn71_58 sn72_58 11.551961
Rsp71_59 sp71_59 sp72_59 11.551961
Rsn71_59 sn71_59 sn72_59 11.551961
Rsp71_60 sp71_60 sp72_60 11.551961
Rsn71_60 sn71_60 sn72_60 11.551961
Rsp71_61 sp71_61 sp72_61 11.551961
Rsn71_61 sn71_61 sn72_61 11.551961
Rsp71_62 sp71_62 sp72_62 11.551961
Rsn71_62 sn71_62 sn72_62 11.551961
Rsp71_63 sp71_63 sp72_63 11.551961
Rsn71_63 sn71_63 sn72_63 11.551961
Rsp71_64 sp71_64 sp72_64 11.551961
Rsn71_64 sn71_64 sn72_64 11.551961
Rsp71_65 sp71_65 sp72_65 11.551961
Rsn71_65 sn71_65 sn72_65 11.551961
Rsp71_66 sp71_66 sp72_66 11.551961
Rsn71_66 sn71_66 sn72_66 11.551961
Rsp71_67 sp71_67 sp72_67 11.551961
Rsn71_67 sn71_67 sn72_67 11.551961
Rsp71_68 sp71_68 sp72_68 11.551961
Rsn71_68 sn71_68 sn72_68 11.551961
Rsp71_69 sp71_69 sp72_69 11.551961
Rsn71_69 sn71_69 sn72_69 11.551961
Rsp71_70 sp71_70 sp72_70 11.551961
Rsn71_70 sn71_70 sn72_70 11.551961
Rsp71_71 sp71_71 sp72_71 11.551961
Rsn71_71 sn71_71 sn72_71 11.551961
Rsp71_72 sp71_72 sp72_72 11.551961
Rsn71_72 sn71_72 sn72_72 11.551961
Rsp71_73 sp71_73 sp72_73 11.551961
Rsn71_73 sn71_73 sn72_73 11.551961
Rsp71_74 sp71_74 sp72_74 11.551961
Rsn71_74 sn71_74 sn72_74 11.551961
Rsp71_75 sp71_75 sp72_75 11.551961
Rsn71_75 sn71_75 sn72_75 11.551961
Rsp71_76 sp71_76 sp72_76 11.551961
Rsn71_76 sn71_76 sn72_76 11.551961
Rsp71_77 sp71_77 sp72_77 11.551961
Rsn71_77 sn71_77 sn72_77 11.551961
Rsp71_78 sp71_78 sp72_78 11.551961
Rsn71_78 sn71_78 sn72_78 11.551961
Rsp71_79 sp71_79 sp72_79 11.551961
Rsn71_79 sn71_79 sn72_79 11.551961
Rsp71_80 sp71_80 sp72_80 11.551961
Rsn71_80 sn71_80 sn72_80 11.551961
Rsp71_81 sp71_81 sp72_81 11.551961
Rsn71_81 sn71_81 sn72_81 11.551961
Rsp71_82 sp71_82 sp72_82 11.551961
Rsn71_82 sn71_82 sn72_82 11.551961
Rsp71_83 sp71_83 sp72_83 11.551961
Rsn71_83 sn71_83 sn72_83 11.551961
Rsp71_84 sp71_84 sp72_84 11.551961
Rsn71_84 sn71_84 sn72_84 11.551961
Rsp72_1 sp72_1 sp73_1 11.551961
Rsn72_1 sn72_1 sn73_1 11.551961
Rsp72_2 sp72_2 sp73_2 11.551961
Rsn72_2 sn72_2 sn73_2 11.551961
Rsp72_3 sp72_3 sp73_3 11.551961
Rsn72_3 sn72_3 sn73_3 11.551961
Rsp72_4 sp72_4 sp73_4 11.551961
Rsn72_4 sn72_4 sn73_4 11.551961
Rsp72_5 sp72_5 sp73_5 11.551961
Rsn72_5 sn72_5 sn73_5 11.551961
Rsp72_6 sp72_6 sp73_6 11.551961
Rsn72_6 sn72_6 sn73_6 11.551961
Rsp72_7 sp72_7 sp73_7 11.551961
Rsn72_7 sn72_7 sn73_7 11.551961
Rsp72_8 sp72_8 sp73_8 11.551961
Rsn72_8 sn72_8 sn73_8 11.551961
Rsp72_9 sp72_9 sp73_9 11.551961
Rsn72_9 sn72_9 sn73_9 11.551961
Rsp72_10 sp72_10 sp73_10 11.551961
Rsn72_10 sn72_10 sn73_10 11.551961
Rsp72_11 sp72_11 sp73_11 11.551961
Rsn72_11 sn72_11 sn73_11 11.551961
Rsp72_12 sp72_12 sp73_12 11.551961
Rsn72_12 sn72_12 sn73_12 11.551961
Rsp72_13 sp72_13 sp73_13 11.551961
Rsn72_13 sn72_13 sn73_13 11.551961
Rsp72_14 sp72_14 sp73_14 11.551961
Rsn72_14 sn72_14 sn73_14 11.551961
Rsp72_15 sp72_15 sp73_15 11.551961
Rsn72_15 sn72_15 sn73_15 11.551961
Rsp72_16 sp72_16 sp73_16 11.551961
Rsn72_16 sn72_16 sn73_16 11.551961
Rsp72_17 sp72_17 sp73_17 11.551961
Rsn72_17 sn72_17 sn73_17 11.551961
Rsp72_18 sp72_18 sp73_18 11.551961
Rsn72_18 sn72_18 sn73_18 11.551961
Rsp72_19 sp72_19 sp73_19 11.551961
Rsn72_19 sn72_19 sn73_19 11.551961
Rsp72_20 sp72_20 sp73_20 11.551961
Rsn72_20 sn72_20 sn73_20 11.551961
Rsp72_21 sp72_21 sp73_21 11.551961
Rsn72_21 sn72_21 sn73_21 11.551961
Rsp72_22 sp72_22 sp73_22 11.551961
Rsn72_22 sn72_22 sn73_22 11.551961
Rsp72_23 sp72_23 sp73_23 11.551961
Rsn72_23 sn72_23 sn73_23 11.551961
Rsp72_24 sp72_24 sp73_24 11.551961
Rsn72_24 sn72_24 sn73_24 11.551961
Rsp72_25 sp72_25 sp73_25 11.551961
Rsn72_25 sn72_25 sn73_25 11.551961
Rsp72_26 sp72_26 sp73_26 11.551961
Rsn72_26 sn72_26 sn73_26 11.551961
Rsp72_27 sp72_27 sp73_27 11.551961
Rsn72_27 sn72_27 sn73_27 11.551961
Rsp72_28 sp72_28 sp73_28 11.551961
Rsn72_28 sn72_28 sn73_28 11.551961
Rsp72_29 sp72_29 sp73_29 11.551961
Rsn72_29 sn72_29 sn73_29 11.551961
Rsp72_30 sp72_30 sp73_30 11.551961
Rsn72_30 sn72_30 sn73_30 11.551961
Rsp72_31 sp72_31 sp73_31 11.551961
Rsn72_31 sn72_31 sn73_31 11.551961
Rsp72_32 sp72_32 sp73_32 11.551961
Rsn72_32 sn72_32 sn73_32 11.551961
Rsp72_33 sp72_33 sp73_33 11.551961
Rsn72_33 sn72_33 sn73_33 11.551961
Rsp72_34 sp72_34 sp73_34 11.551961
Rsn72_34 sn72_34 sn73_34 11.551961
Rsp72_35 sp72_35 sp73_35 11.551961
Rsn72_35 sn72_35 sn73_35 11.551961
Rsp72_36 sp72_36 sp73_36 11.551961
Rsn72_36 sn72_36 sn73_36 11.551961
Rsp72_37 sp72_37 sp73_37 11.551961
Rsn72_37 sn72_37 sn73_37 11.551961
Rsp72_38 sp72_38 sp73_38 11.551961
Rsn72_38 sn72_38 sn73_38 11.551961
Rsp72_39 sp72_39 sp73_39 11.551961
Rsn72_39 sn72_39 sn73_39 11.551961
Rsp72_40 sp72_40 sp73_40 11.551961
Rsn72_40 sn72_40 sn73_40 11.551961
Rsp72_41 sp72_41 sp73_41 11.551961
Rsn72_41 sn72_41 sn73_41 11.551961
Rsp72_42 sp72_42 sp73_42 11.551961
Rsn72_42 sn72_42 sn73_42 11.551961
Rsp72_43 sp72_43 sp73_43 11.551961
Rsn72_43 sn72_43 sn73_43 11.551961
Rsp72_44 sp72_44 sp73_44 11.551961
Rsn72_44 sn72_44 sn73_44 11.551961
Rsp72_45 sp72_45 sp73_45 11.551961
Rsn72_45 sn72_45 sn73_45 11.551961
Rsp72_46 sp72_46 sp73_46 11.551961
Rsn72_46 sn72_46 sn73_46 11.551961
Rsp72_47 sp72_47 sp73_47 11.551961
Rsn72_47 sn72_47 sn73_47 11.551961
Rsp72_48 sp72_48 sp73_48 11.551961
Rsn72_48 sn72_48 sn73_48 11.551961
Rsp72_49 sp72_49 sp73_49 11.551961
Rsn72_49 sn72_49 sn73_49 11.551961
Rsp72_50 sp72_50 sp73_50 11.551961
Rsn72_50 sn72_50 sn73_50 11.551961
Rsp72_51 sp72_51 sp73_51 11.551961
Rsn72_51 sn72_51 sn73_51 11.551961
Rsp72_52 sp72_52 sp73_52 11.551961
Rsn72_52 sn72_52 sn73_52 11.551961
Rsp72_53 sp72_53 sp73_53 11.551961
Rsn72_53 sn72_53 sn73_53 11.551961
Rsp72_54 sp72_54 sp73_54 11.551961
Rsn72_54 sn72_54 sn73_54 11.551961
Rsp72_55 sp72_55 sp73_55 11.551961
Rsn72_55 sn72_55 sn73_55 11.551961
Rsp72_56 sp72_56 sp73_56 11.551961
Rsn72_56 sn72_56 sn73_56 11.551961
Rsp72_57 sp72_57 sp73_57 11.551961
Rsn72_57 sn72_57 sn73_57 11.551961
Rsp72_58 sp72_58 sp73_58 11.551961
Rsn72_58 sn72_58 sn73_58 11.551961
Rsp72_59 sp72_59 sp73_59 11.551961
Rsn72_59 sn72_59 sn73_59 11.551961
Rsp72_60 sp72_60 sp73_60 11.551961
Rsn72_60 sn72_60 sn73_60 11.551961
Rsp72_61 sp72_61 sp73_61 11.551961
Rsn72_61 sn72_61 sn73_61 11.551961
Rsp72_62 sp72_62 sp73_62 11.551961
Rsn72_62 sn72_62 sn73_62 11.551961
Rsp72_63 sp72_63 sp73_63 11.551961
Rsn72_63 sn72_63 sn73_63 11.551961
Rsp72_64 sp72_64 sp73_64 11.551961
Rsn72_64 sn72_64 sn73_64 11.551961
Rsp72_65 sp72_65 sp73_65 11.551961
Rsn72_65 sn72_65 sn73_65 11.551961
Rsp72_66 sp72_66 sp73_66 11.551961
Rsn72_66 sn72_66 sn73_66 11.551961
Rsp72_67 sp72_67 sp73_67 11.551961
Rsn72_67 sn72_67 sn73_67 11.551961
Rsp72_68 sp72_68 sp73_68 11.551961
Rsn72_68 sn72_68 sn73_68 11.551961
Rsp72_69 sp72_69 sp73_69 11.551961
Rsn72_69 sn72_69 sn73_69 11.551961
Rsp72_70 sp72_70 sp73_70 11.551961
Rsn72_70 sn72_70 sn73_70 11.551961
Rsp72_71 sp72_71 sp73_71 11.551961
Rsn72_71 sn72_71 sn73_71 11.551961
Rsp72_72 sp72_72 sp73_72 11.551961
Rsn72_72 sn72_72 sn73_72 11.551961
Rsp72_73 sp72_73 sp73_73 11.551961
Rsn72_73 sn72_73 sn73_73 11.551961
Rsp72_74 sp72_74 sp73_74 11.551961
Rsn72_74 sn72_74 sn73_74 11.551961
Rsp72_75 sp72_75 sp73_75 11.551961
Rsn72_75 sn72_75 sn73_75 11.551961
Rsp72_76 sp72_76 sp73_76 11.551961
Rsn72_76 sn72_76 sn73_76 11.551961
Rsp72_77 sp72_77 sp73_77 11.551961
Rsn72_77 sn72_77 sn73_77 11.551961
Rsp72_78 sp72_78 sp73_78 11.551961
Rsn72_78 sn72_78 sn73_78 11.551961
Rsp72_79 sp72_79 sp73_79 11.551961
Rsn72_79 sn72_79 sn73_79 11.551961
Rsp72_80 sp72_80 sp73_80 11.551961
Rsn72_80 sn72_80 sn73_80 11.551961
Rsp72_81 sp72_81 sp73_81 11.551961
Rsn72_81 sn72_81 sn73_81 11.551961
Rsp72_82 sp72_82 sp73_82 11.551961
Rsn72_82 sn72_82 sn73_82 11.551961
Rsp72_83 sp72_83 sp73_83 11.551961
Rsn72_83 sn72_83 sn73_83 11.551961
Rsp72_84 sp72_84 sp73_84 11.551961
Rsn72_84 sn72_84 sn73_84 11.551961
Rsp73_1 sp73_1 sp74_1 11.551961
Rsn73_1 sn73_1 sn74_1 11.551961
Rsp73_2 sp73_2 sp74_2 11.551961
Rsn73_2 sn73_2 sn74_2 11.551961
Rsp73_3 sp73_3 sp74_3 11.551961
Rsn73_3 sn73_3 sn74_3 11.551961
Rsp73_4 sp73_4 sp74_4 11.551961
Rsn73_4 sn73_4 sn74_4 11.551961
Rsp73_5 sp73_5 sp74_5 11.551961
Rsn73_5 sn73_5 sn74_5 11.551961
Rsp73_6 sp73_6 sp74_6 11.551961
Rsn73_6 sn73_6 sn74_6 11.551961
Rsp73_7 sp73_7 sp74_7 11.551961
Rsn73_7 sn73_7 sn74_7 11.551961
Rsp73_8 sp73_8 sp74_8 11.551961
Rsn73_8 sn73_8 sn74_8 11.551961
Rsp73_9 sp73_9 sp74_9 11.551961
Rsn73_9 sn73_9 sn74_9 11.551961
Rsp73_10 sp73_10 sp74_10 11.551961
Rsn73_10 sn73_10 sn74_10 11.551961
Rsp73_11 sp73_11 sp74_11 11.551961
Rsn73_11 sn73_11 sn74_11 11.551961
Rsp73_12 sp73_12 sp74_12 11.551961
Rsn73_12 sn73_12 sn74_12 11.551961
Rsp73_13 sp73_13 sp74_13 11.551961
Rsn73_13 sn73_13 sn74_13 11.551961
Rsp73_14 sp73_14 sp74_14 11.551961
Rsn73_14 sn73_14 sn74_14 11.551961
Rsp73_15 sp73_15 sp74_15 11.551961
Rsn73_15 sn73_15 sn74_15 11.551961
Rsp73_16 sp73_16 sp74_16 11.551961
Rsn73_16 sn73_16 sn74_16 11.551961
Rsp73_17 sp73_17 sp74_17 11.551961
Rsn73_17 sn73_17 sn74_17 11.551961
Rsp73_18 sp73_18 sp74_18 11.551961
Rsn73_18 sn73_18 sn74_18 11.551961
Rsp73_19 sp73_19 sp74_19 11.551961
Rsn73_19 sn73_19 sn74_19 11.551961
Rsp73_20 sp73_20 sp74_20 11.551961
Rsn73_20 sn73_20 sn74_20 11.551961
Rsp73_21 sp73_21 sp74_21 11.551961
Rsn73_21 sn73_21 sn74_21 11.551961
Rsp73_22 sp73_22 sp74_22 11.551961
Rsn73_22 sn73_22 sn74_22 11.551961
Rsp73_23 sp73_23 sp74_23 11.551961
Rsn73_23 sn73_23 sn74_23 11.551961
Rsp73_24 sp73_24 sp74_24 11.551961
Rsn73_24 sn73_24 sn74_24 11.551961
Rsp73_25 sp73_25 sp74_25 11.551961
Rsn73_25 sn73_25 sn74_25 11.551961
Rsp73_26 sp73_26 sp74_26 11.551961
Rsn73_26 sn73_26 sn74_26 11.551961
Rsp73_27 sp73_27 sp74_27 11.551961
Rsn73_27 sn73_27 sn74_27 11.551961
Rsp73_28 sp73_28 sp74_28 11.551961
Rsn73_28 sn73_28 sn74_28 11.551961
Rsp73_29 sp73_29 sp74_29 11.551961
Rsn73_29 sn73_29 sn74_29 11.551961
Rsp73_30 sp73_30 sp74_30 11.551961
Rsn73_30 sn73_30 sn74_30 11.551961
Rsp73_31 sp73_31 sp74_31 11.551961
Rsn73_31 sn73_31 sn74_31 11.551961
Rsp73_32 sp73_32 sp74_32 11.551961
Rsn73_32 sn73_32 sn74_32 11.551961
Rsp73_33 sp73_33 sp74_33 11.551961
Rsn73_33 sn73_33 sn74_33 11.551961
Rsp73_34 sp73_34 sp74_34 11.551961
Rsn73_34 sn73_34 sn74_34 11.551961
Rsp73_35 sp73_35 sp74_35 11.551961
Rsn73_35 sn73_35 sn74_35 11.551961
Rsp73_36 sp73_36 sp74_36 11.551961
Rsn73_36 sn73_36 sn74_36 11.551961
Rsp73_37 sp73_37 sp74_37 11.551961
Rsn73_37 sn73_37 sn74_37 11.551961
Rsp73_38 sp73_38 sp74_38 11.551961
Rsn73_38 sn73_38 sn74_38 11.551961
Rsp73_39 sp73_39 sp74_39 11.551961
Rsn73_39 sn73_39 sn74_39 11.551961
Rsp73_40 sp73_40 sp74_40 11.551961
Rsn73_40 sn73_40 sn74_40 11.551961
Rsp73_41 sp73_41 sp74_41 11.551961
Rsn73_41 sn73_41 sn74_41 11.551961
Rsp73_42 sp73_42 sp74_42 11.551961
Rsn73_42 sn73_42 sn74_42 11.551961
Rsp73_43 sp73_43 sp74_43 11.551961
Rsn73_43 sn73_43 sn74_43 11.551961
Rsp73_44 sp73_44 sp74_44 11.551961
Rsn73_44 sn73_44 sn74_44 11.551961
Rsp73_45 sp73_45 sp74_45 11.551961
Rsn73_45 sn73_45 sn74_45 11.551961
Rsp73_46 sp73_46 sp74_46 11.551961
Rsn73_46 sn73_46 sn74_46 11.551961
Rsp73_47 sp73_47 sp74_47 11.551961
Rsn73_47 sn73_47 sn74_47 11.551961
Rsp73_48 sp73_48 sp74_48 11.551961
Rsn73_48 sn73_48 sn74_48 11.551961
Rsp73_49 sp73_49 sp74_49 11.551961
Rsn73_49 sn73_49 sn74_49 11.551961
Rsp73_50 sp73_50 sp74_50 11.551961
Rsn73_50 sn73_50 sn74_50 11.551961
Rsp73_51 sp73_51 sp74_51 11.551961
Rsn73_51 sn73_51 sn74_51 11.551961
Rsp73_52 sp73_52 sp74_52 11.551961
Rsn73_52 sn73_52 sn74_52 11.551961
Rsp73_53 sp73_53 sp74_53 11.551961
Rsn73_53 sn73_53 sn74_53 11.551961
Rsp73_54 sp73_54 sp74_54 11.551961
Rsn73_54 sn73_54 sn74_54 11.551961
Rsp73_55 sp73_55 sp74_55 11.551961
Rsn73_55 sn73_55 sn74_55 11.551961
Rsp73_56 sp73_56 sp74_56 11.551961
Rsn73_56 sn73_56 sn74_56 11.551961
Rsp73_57 sp73_57 sp74_57 11.551961
Rsn73_57 sn73_57 sn74_57 11.551961
Rsp73_58 sp73_58 sp74_58 11.551961
Rsn73_58 sn73_58 sn74_58 11.551961
Rsp73_59 sp73_59 sp74_59 11.551961
Rsn73_59 sn73_59 sn74_59 11.551961
Rsp73_60 sp73_60 sp74_60 11.551961
Rsn73_60 sn73_60 sn74_60 11.551961
Rsp73_61 sp73_61 sp74_61 11.551961
Rsn73_61 sn73_61 sn74_61 11.551961
Rsp73_62 sp73_62 sp74_62 11.551961
Rsn73_62 sn73_62 sn74_62 11.551961
Rsp73_63 sp73_63 sp74_63 11.551961
Rsn73_63 sn73_63 sn74_63 11.551961
Rsp73_64 sp73_64 sp74_64 11.551961
Rsn73_64 sn73_64 sn74_64 11.551961
Rsp73_65 sp73_65 sp74_65 11.551961
Rsn73_65 sn73_65 sn74_65 11.551961
Rsp73_66 sp73_66 sp74_66 11.551961
Rsn73_66 sn73_66 sn74_66 11.551961
Rsp73_67 sp73_67 sp74_67 11.551961
Rsn73_67 sn73_67 sn74_67 11.551961
Rsp73_68 sp73_68 sp74_68 11.551961
Rsn73_68 sn73_68 sn74_68 11.551961
Rsp73_69 sp73_69 sp74_69 11.551961
Rsn73_69 sn73_69 sn74_69 11.551961
Rsp73_70 sp73_70 sp74_70 11.551961
Rsn73_70 sn73_70 sn74_70 11.551961
Rsp73_71 sp73_71 sp74_71 11.551961
Rsn73_71 sn73_71 sn74_71 11.551961
Rsp73_72 sp73_72 sp74_72 11.551961
Rsn73_72 sn73_72 sn74_72 11.551961
Rsp73_73 sp73_73 sp74_73 11.551961
Rsn73_73 sn73_73 sn74_73 11.551961
Rsp73_74 sp73_74 sp74_74 11.551961
Rsn73_74 sn73_74 sn74_74 11.551961
Rsp73_75 sp73_75 sp74_75 11.551961
Rsn73_75 sn73_75 sn74_75 11.551961
Rsp73_76 sp73_76 sp74_76 11.551961
Rsn73_76 sn73_76 sn74_76 11.551961
Rsp73_77 sp73_77 sp74_77 11.551961
Rsn73_77 sn73_77 sn74_77 11.551961
Rsp73_78 sp73_78 sp74_78 11.551961
Rsn73_78 sn73_78 sn74_78 11.551961
Rsp73_79 sp73_79 sp74_79 11.551961
Rsn73_79 sn73_79 sn74_79 11.551961
Rsp73_80 sp73_80 sp74_80 11.551961
Rsn73_80 sn73_80 sn74_80 11.551961
Rsp73_81 sp73_81 sp74_81 11.551961
Rsn73_81 sn73_81 sn74_81 11.551961
Rsp73_82 sp73_82 sp74_82 11.551961
Rsn73_82 sn73_82 sn74_82 11.551961
Rsp73_83 sp73_83 sp74_83 11.551961
Rsn73_83 sn73_83 sn74_83 11.551961
Rsp73_84 sp73_84 sp74_84 11.551961
Rsn73_84 sn73_84 sn74_84 11.551961
Rsp74_1 sp74_1 sp75_1 11.551961
Rsn74_1 sn74_1 sn75_1 11.551961
Rsp74_2 sp74_2 sp75_2 11.551961
Rsn74_2 sn74_2 sn75_2 11.551961
Rsp74_3 sp74_3 sp75_3 11.551961
Rsn74_3 sn74_3 sn75_3 11.551961
Rsp74_4 sp74_4 sp75_4 11.551961
Rsn74_4 sn74_4 sn75_4 11.551961
Rsp74_5 sp74_5 sp75_5 11.551961
Rsn74_5 sn74_5 sn75_5 11.551961
Rsp74_6 sp74_6 sp75_6 11.551961
Rsn74_6 sn74_6 sn75_6 11.551961
Rsp74_7 sp74_7 sp75_7 11.551961
Rsn74_7 sn74_7 sn75_7 11.551961
Rsp74_8 sp74_8 sp75_8 11.551961
Rsn74_8 sn74_8 sn75_8 11.551961
Rsp74_9 sp74_9 sp75_9 11.551961
Rsn74_9 sn74_9 sn75_9 11.551961
Rsp74_10 sp74_10 sp75_10 11.551961
Rsn74_10 sn74_10 sn75_10 11.551961
Rsp74_11 sp74_11 sp75_11 11.551961
Rsn74_11 sn74_11 sn75_11 11.551961
Rsp74_12 sp74_12 sp75_12 11.551961
Rsn74_12 sn74_12 sn75_12 11.551961
Rsp74_13 sp74_13 sp75_13 11.551961
Rsn74_13 sn74_13 sn75_13 11.551961
Rsp74_14 sp74_14 sp75_14 11.551961
Rsn74_14 sn74_14 sn75_14 11.551961
Rsp74_15 sp74_15 sp75_15 11.551961
Rsn74_15 sn74_15 sn75_15 11.551961
Rsp74_16 sp74_16 sp75_16 11.551961
Rsn74_16 sn74_16 sn75_16 11.551961
Rsp74_17 sp74_17 sp75_17 11.551961
Rsn74_17 sn74_17 sn75_17 11.551961
Rsp74_18 sp74_18 sp75_18 11.551961
Rsn74_18 sn74_18 sn75_18 11.551961
Rsp74_19 sp74_19 sp75_19 11.551961
Rsn74_19 sn74_19 sn75_19 11.551961
Rsp74_20 sp74_20 sp75_20 11.551961
Rsn74_20 sn74_20 sn75_20 11.551961
Rsp74_21 sp74_21 sp75_21 11.551961
Rsn74_21 sn74_21 sn75_21 11.551961
Rsp74_22 sp74_22 sp75_22 11.551961
Rsn74_22 sn74_22 sn75_22 11.551961
Rsp74_23 sp74_23 sp75_23 11.551961
Rsn74_23 sn74_23 sn75_23 11.551961
Rsp74_24 sp74_24 sp75_24 11.551961
Rsn74_24 sn74_24 sn75_24 11.551961
Rsp74_25 sp74_25 sp75_25 11.551961
Rsn74_25 sn74_25 sn75_25 11.551961
Rsp74_26 sp74_26 sp75_26 11.551961
Rsn74_26 sn74_26 sn75_26 11.551961
Rsp74_27 sp74_27 sp75_27 11.551961
Rsn74_27 sn74_27 sn75_27 11.551961
Rsp74_28 sp74_28 sp75_28 11.551961
Rsn74_28 sn74_28 sn75_28 11.551961
Rsp74_29 sp74_29 sp75_29 11.551961
Rsn74_29 sn74_29 sn75_29 11.551961
Rsp74_30 sp74_30 sp75_30 11.551961
Rsn74_30 sn74_30 sn75_30 11.551961
Rsp74_31 sp74_31 sp75_31 11.551961
Rsn74_31 sn74_31 sn75_31 11.551961
Rsp74_32 sp74_32 sp75_32 11.551961
Rsn74_32 sn74_32 sn75_32 11.551961
Rsp74_33 sp74_33 sp75_33 11.551961
Rsn74_33 sn74_33 sn75_33 11.551961
Rsp74_34 sp74_34 sp75_34 11.551961
Rsn74_34 sn74_34 sn75_34 11.551961
Rsp74_35 sp74_35 sp75_35 11.551961
Rsn74_35 sn74_35 sn75_35 11.551961
Rsp74_36 sp74_36 sp75_36 11.551961
Rsn74_36 sn74_36 sn75_36 11.551961
Rsp74_37 sp74_37 sp75_37 11.551961
Rsn74_37 sn74_37 sn75_37 11.551961
Rsp74_38 sp74_38 sp75_38 11.551961
Rsn74_38 sn74_38 sn75_38 11.551961
Rsp74_39 sp74_39 sp75_39 11.551961
Rsn74_39 sn74_39 sn75_39 11.551961
Rsp74_40 sp74_40 sp75_40 11.551961
Rsn74_40 sn74_40 sn75_40 11.551961
Rsp74_41 sp74_41 sp75_41 11.551961
Rsn74_41 sn74_41 sn75_41 11.551961
Rsp74_42 sp74_42 sp75_42 11.551961
Rsn74_42 sn74_42 sn75_42 11.551961
Rsp74_43 sp74_43 sp75_43 11.551961
Rsn74_43 sn74_43 sn75_43 11.551961
Rsp74_44 sp74_44 sp75_44 11.551961
Rsn74_44 sn74_44 sn75_44 11.551961
Rsp74_45 sp74_45 sp75_45 11.551961
Rsn74_45 sn74_45 sn75_45 11.551961
Rsp74_46 sp74_46 sp75_46 11.551961
Rsn74_46 sn74_46 sn75_46 11.551961
Rsp74_47 sp74_47 sp75_47 11.551961
Rsn74_47 sn74_47 sn75_47 11.551961
Rsp74_48 sp74_48 sp75_48 11.551961
Rsn74_48 sn74_48 sn75_48 11.551961
Rsp74_49 sp74_49 sp75_49 11.551961
Rsn74_49 sn74_49 sn75_49 11.551961
Rsp74_50 sp74_50 sp75_50 11.551961
Rsn74_50 sn74_50 sn75_50 11.551961
Rsp74_51 sp74_51 sp75_51 11.551961
Rsn74_51 sn74_51 sn75_51 11.551961
Rsp74_52 sp74_52 sp75_52 11.551961
Rsn74_52 sn74_52 sn75_52 11.551961
Rsp74_53 sp74_53 sp75_53 11.551961
Rsn74_53 sn74_53 sn75_53 11.551961
Rsp74_54 sp74_54 sp75_54 11.551961
Rsn74_54 sn74_54 sn75_54 11.551961
Rsp74_55 sp74_55 sp75_55 11.551961
Rsn74_55 sn74_55 sn75_55 11.551961
Rsp74_56 sp74_56 sp75_56 11.551961
Rsn74_56 sn74_56 sn75_56 11.551961
Rsp74_57 sp74_57 sp75_57 11.551961
Rsn74_57 sn74_57 sn75_57 11.551961
Rsp74_58 sp74_58 sp75_58 11.551961
Rsn74_58 sn74_58 sn75_58 11.551961
Rsp74_59 sp74_59 sp75_59 11.551961
Rsn74_59 sn74_59 sn75_59 11.551961
Rsp74_60 sp74_60 sp75_60 11.551961
Rsn74_60 sn74_60 sn75_60 11.551961
Rsp74_61 sp74_61 sp75_61 11.551961
Rsn74_61 sn74_61 sn75_61 11.551961
Rsp74_62 sp74_62 sp75_62 11.551961
Rsn74_62 sn74_62 sn75_62 11.551961
Rsp74_63 sp74_63 sp75_63 11.551961
Rsn74_63 sn74_63 sn75_63 11.551961
Rsp74_64 sp74_64 sp75_64 11.551961
Rsn74_64 sn74_64 sn75_64 11.551961
Rsp74_65 sp74_65 sp75_65 11.551961
Rsn74_65 sn74_65 sn75_65 11.551961
Rsp74_66 sp74_66 sp75_66 11.551961
Rsn74_66 sn74_66 sn75_66 11.551961
Rsp74_67 sp74_67 sp75_67 11.551961
Rsn74_67 sn74_67 sn75_67 11.551961
Rsp74_68 sp74_68 sp75_68 11.551961
Rsn74_68 sn74_68 sn75_68 11.551961
Rsp74_69 sp74_69 sp75_69 11.551961
Rsn74_69 sn74_69 sn75_69 11.551961
Rsp74_70 sp74_70 sp75_70 11.551961
Rsn74_70 sn74_70 sn75_70 11.551961
Rsp74_71 sp74_71 sp75_71 11.551961
Rsn74_71 sn74_71 sn75_71 11.551961
Rsp74_72 sp74_72 sp75_72 11.551961
Rsn74_72 sn74_72 sn75_72 11.551961
Rsp74_73 sp74_73 sp75_73 11.551961
Rsn74_73 sn74_73 sn75_73 11.551961
Rsp74_74 sp74_74 sp75_74 11.551961
Rsn74_74 sn74_74 sn75_74 11.551961
Rsp74_75 sp74_75 sp75_75 11.551961
Rsn74_75 sn74_75 sn75_75 11.551961
Rsp74_76 sp74_76 sp75_76 11.551961
Rsn74_76 sn74_76 sn75_76 11.551961
Rsp74_77 sp74_77 sp75_77 11.551961
Rsn74_77 sn74_77 sn75_77 11.551961
Rsp74_78 sp74_78 sp75_78 11.551961
Rsn74_78 sn74_78 sn75_78 11.551961
Rsp74_79 sp74_79 sp75_79 11.551961
Rsn74_79 sn74_79 sn75_79 11.551961
Rsp74_80 sp74_80 sp75_80 11.551961
Rsn74_80 sn74_80 sn75_80 11.551961
Rsp74_81 sp74_81 sp75_81 11.551961
Rsn74_81 sn74_81 sn75_81 11.551961
Rsp74_82 sp74_82 sp75_82 11.551961
Rsn74_82 sn74_82 sn75_82 11.551961
Rsp74_83 sp74_83 sp75_83 11.551961
Rsn74_83 sn74_83 sn75_83 11.551961
Rsp74_84 sp74_84 sp75_84 11.551961
Rsn74_84 sn74_84 sn75_84 11.551961
Rsp75_1 sp75_1 sp76_1 11.551961
Rsn75_1 sn75_1 sn76_1 11.551961
Rsp75_2 sp75_2 sp76_2 11.551961
Rsn75_2 sn75_2 sn76_2 11.551961
Rsp75_3 sp75_3 sp76_3 11.551961
Rsn75_3 sn75_3 sn76_3 11.551961
Rsp75_4 sp75_4 sp76_4 11.551961
Rsn75_4 sn75_4 sn76_4 11.551961
Rsp75_5 sp75_5 sp76_5 11.551961
Rsn75_5 sn75_5 sn76_5 11.551961
Rsp75_6 sp75_6 sp76_6 11.551961
Rsn75_6 sn75_6 sn76_6 11.551961
Rsp75_7 sp75_7 sp76_7 11.551961
Rsn75_7 sn75_7 sn76_7 11.551961
Rsp75_8 sp75_8 sp76_8 11.551961
Rsn75_8 sn75_8 sn76_8 11.551961
Rsp75_9 sp75_9 sp76_9 11.551961
Rsn75_9 sn75_9 sn76_9 11.551961
Rsp75_10 sp75_10 sp76_10 11.551961
Rsn75_10 sn75_10 sn76_10 11.551961
Rsp75_11 sp75_11 sp76_11 11.551961
Rsn75_11 sn75_11 sn76_11 11.551961
Rsp75_12 sp75_12 sp76_12 11.551961
Rsn75_12 sn75_12 sn76_12 11.551961
Rsp75_13 sp75_13 sp76_13 11.551961
Rsn75_13 sn75_13 sn76_13 11.551961
Rsp75_14 sp75_14 sp76_14 11.551961
Rsn75_14 sn75_14 sn76_14 11.551961
Rsp75_15 sp75_15 sp76_15 11.551961
Rsn75_15 sn75_15 sn76_15 11.551961
Rsp75_16 sp75_16 sp76_16 11.551961
Rsn75_16 sn75_16 sn76_16 11.551961
Rsp75_17 sp75_17 sp76_17 11.551961
Rsn75_17 sn75_17 sn76_17 11.551961
Rsp75_18 sp75_18 sp76_18 11.551961
Rsn75_18 sn75_18 sn76_18 11.551961
Rsp75_19 sp75_19 sp76_19 11.551961
Rsn75_19 sn75_19 sn76_19 11.551961
Rsp75_20 sp75_20 sp76_20 11.551961
Rsn75_20 sn75_20 sn76_20 11.551961
Rsp75_21 sp75_21 sp76_21 11.551961
Rsn75_21 sn75_21 sn76_21 11.551961
Rsp75_22 sp75_22 sp76_22 11.551961
Rsn75_22 sn75_22 sn76_22 11.551961
Rsp75_23 sp75_23 sp76_23 11.551961
Rsn75_23 sn75_23 sn76_23 11.551961
Rsp75_24 sp75_24 sp76_24 11.551961
Rsn75_24 sn75_24 sn76_24 11.551961
Rsp75_25 sp75_25 sp76_25 11.551961
Rsn75_25 sn75_25 sn76_25 11.551961
Rsp75_26 sp75_26 sp76_26 11.551961
Rsn75_26 sn75_26 sn76_26 11.551961
Rsp75_27 sp75_27 sp76_27 11.551961
Rsn75_27 sn75_27 sn76_27 11.551961
Rsp75_28 sp75_28 sp76_28 11.551961
Rsn75_28 sn75_28 sn76_28 11.551961
Rsp75_29 sp75_29 sp76_29 11.551961
Rsn75_29 sn75_29 sn76_29 11.551961
Rsp75_30 sp75_30 sp76_30 11.551961
Rsn75_30 sn75_30 sn76_30 11.551961
Rsp75_31 sp75_31 sp76_31 11.551961
Rsn75_31 sn75_31 sn76_31 11.551961
Rsp75_32 sp75_32 sp76_32 11.551961
Rsn75_32 sn75_32 sn76_32 11.551961
Rsp75_33 sp75_33 sp76_33 11.551961
Rsn75_33 sn75_33 sn76_33 11.551961
Rsp75_34 sp75_34 sp76_34 11.551961
Rsn75_34 sn75_34 sn76_34 11.551961
Rsp75_35 sp75_35 sp76_35 11.551961
Rsn75_35 sn75_35 sn76_35 11.551961
Rsp75_36 sp75_36 sp76_36 11.551961
Rsn75_36 sn75_36 sn76_36 11.551961
Rsp75_37 sp75_37 sp76_37 11.551961
Rsn75_37 sn75_37 sn76_37 11.551961
Rsp75_38 sp75_38 sp76_38 11.551961
Rsn75_38 sn75_38 sn76_38 11.551961
Rsp75_39 sp75_39 sp76_39 11.551961
Rsn75_39 sn75_39 sn76_39 11.551961
Rsp75_40 sp75_40 sp76_40 11.551961
Rsn75_40 sn75_40 sn76_40 11.551961
Rsp75_41 sp75_41 sp76_41 11.551961
Rsn75_41 sn75_41 sn76_41 11.551961
Rsp75_42 sp75_42 sp76_42 11.551961
Rsn75_42 sn75_42 sn76_42 11.551961
Rsp75_43 sp75_43 sp76_43 11.551961
Rsn75_43 sn75_43 sn76_43 11.551961
Rsp75_44 sp75_44 sp76_44 11.551961
Rsn75_44 sn75_44 sn76_44 11.551961
Rsp75_45 sp75_45 sp76_45 11.551961
Rsn75_45 sn75_45 sn76_45 11.551961
Rsp75_46 sp75_46 sp76_46 11.551961
Rsn75_46 sn75_46 sn76_46 11.551961
Rsp75_47 sp75_47 sp76_47 11.551961
Rsn75_47 sn75_47 sn76_47 11.551961
Rsp75_48 sp75_48 sp76_48 11.551961
Rsn75_48 sn75_48 sn76_48 11.551961
Rsp75_49 sp75_49 sp76_49 11.551961
Rsn75_49 sn75_49 sn76_49 11.551961
Rsp75_50 sp75_50 sp76_50 11.551961
Rsn75_50 sn75_50 sn76_50 11.551961
Rsp75_51 sp75_51 sp76_51 11.551961
Rsn75_51 sn75_51 sn76_51 11.551961
Rsp75_52 sp75_52 sp76_52 11.551961
Rsn75_52 sn75_52 sn76_52 11.551961
Rsp75_53 sp75_53 sp76_53 11.551961
Rsn75_53 sn75_53 sn76_53 11.551961
Rsp75_54 sp75_54 sp76_54 11.551961
Rsn75_54 sn75_54 sn76_54 11.551961
Rsp75_55 sp75_55 sp76_55 11.551961
Rsn75_55 sn75_55 sn76_55 11.551961
Rsp75_56 sp75_56 sp76_56 11.551961
Rsn75_56 sn75_56 sn76_56 11.551961
Rsp75_57 sp75_57 sp76_57 11.551961
Rsn75_57 sn75_57 sn76_57 11.551961
Rsp75_58 sp75_58 sp76_58 11.551961
Rsn75_58 sn75_58 sn76_58 11.551961
Rsp75_59 sp75_59 sp76_59 11.551961
Rsn75_59 sn75_59 sn76_59 11.551961
Rsp75_60 sp75_60 sp76_60 11.551961
Rsn75_60 sn75_60 sn76_60 11.551961
Rsp75_61 sp75_61 sp76_61 11.551961
Rsn75_61 sn75_61 sn76_61 11.551961
Rsp75_62 sp75_62 sp76_62 11.551961
Rsn75_62 sn75_62 sn76_62 11.551961
Rsp75_63 sp75_63 sp76_63 11.551961
Rsn75_63 sn75_63 sn76_63 11.551961
Rsp75_64 sp75_64 sp76_64 11.551961
Rsn75_64 sn75_64 sn76_64 11.551961
Rsp75_65 sp75_65 sp76_65 11.551961
Rsn75_65 sn75_65 sn76_65 11.551961
Rsp75_66 sp75_66 sp76_66 11.551961
Rsn75_66 sn75_66 sn76_66 11.551961
Rsp75_67 sp75_67 sp76_67 11.551961
Rsn75_67 sn75_67 sn76_67 11.551961
Rsp75_68 sp75_68 sp76_68 11.551961
Rsn75_68 sn75_68 sn76_68 11.551961
Rsp75_69 sp75_69 sp76_69 11.551961
Rsn75_69 sn75_69 sn76_69 11.551961
Rsp75_70 sp75_70 sp76_70 11.551961
Rsn75_70 sn75_70 sn76_70 11.551961
Rsp75_71 sp75_71 sp76_71 11.551961
Rsn75_71 sn75_71 sn76_71 11.551961
Rsp75_72 sp75_72 sp76_72 11.551961
Rsn75_72 sn75_72 sn76_72 11.551961
Rsp75_73 sp75_73 sp76_73 11.551961
Rsn75_73 sn75_73 sn76_73 11.551961
Rsp75_74 sp75_74 sp76_74 11.551961
Rsn75_74 sn75_74 sn76_74 11.551961
Rsp75_75 sp75_75 sp76_75 11.551961
Rsn75_75 sn75_75 sn76_75 11.551961
Rsp75_76 sp75_76 sp76_76 11.551961
Rsn75_76 sn75_76 sn76_76 11.551961
Rsp75_77 sp75_77 sp76_77 11.551961
Rsn75_77 sn75_77 sn76_77 11.551961
Rsp75_78 sp75_78 sp76_78 11.551961
Rsn75_78 sn75_78 sn76_78 11.551961
Rsp75_79 sp75_79 sp76_79 11.551961
Rsn75_79 sn75_79 sn76_79 11.551961
Rsp75_80 sp75_80 sp76_80 11.551961
Rsn75_80 sn75_80 sn76_80 11.551961
Rsp75_81 sp75_81 sp76_81 11.551961
Rsn75_81 sn75_81 sn76_81 11.551961
Rsp75_82 sp75_82 sp76_82 11.551961
Rsn75_82 sn75_82 sn76_82 11.551961
Rsp75_83 sp75_83 sp76_83 11.551961
Rsn75_83 sn75_83 sn76_83 11.551961
Rsp75_84 sp75_84 sp76_84 11.551961
Rsn75_84 sn75_84 sn76_84 11.551961
Rsp76_1 sp76_1 sp77_1 11.551961
Rsn76_1 sn76_1 sn77_1 11.551961
Rsp76_2 sp76_2 sp77_2 11.551961
Rsn76_2 sn76_2 sn77_2 11.551961
Rsp76_3 sp76_3 sp77_3 11.551961
Rsn76_3 sn76_3 sn77_3 11.551961
Rsp76_4 sp76_4 sp77_4 11.551961
Rsn76_4 sn76_4 sn77_4 11.551961
Rsp76_5 sp76_5 sp77_5 11.551961
Rsn76_5 sn76_5 sn77_5 11.551961
Rsp76_6 sp76_6 sp77_6 11.551961
Rsn76_6 sn76_6 sn77_6 11.551961
Rsp76_7 sp76_7 sp77_7 11.551961
Rsn76_7 sn76_7 sn77_7 11.551961
Rsp76_8 sp76_8 sp77_8 11.551961
Rsn76_8 sn76_8 sn77_8 11.551961
Rsp76_9 sp76_9 sp77_9 11.551961
Rsn76_9 sn76_9 sn77_9 11.551961
Rsp76_10 sp76_10 sp77_10 11.551961
Rsn76_10 sn76_10 sn77_10 11.551961
Rsp76_11 sp76_11 sp77_11 11.551961
Rsn76_11 sn76_11 sn77_11 11.551961
Rsp76_12 sp76_12 sp77_12 11.551961
Rsn76_12 sn76_12 sn77_12 11.551961
Rsp76_13 sp76_13 sp77_13 11.551961
Rsn76_13 sn76_13 sn77_13 11.551961
Rsp76_14 sp76_14 sp77_14 11.551961
Rsn76_14 sn76_14 sn77_14 11.551961
Rsp76_15 sp76_15 sp77_15 11.551961
Rsn76_15 sn76_15 sn77_15 11.551961
Rsp76_16 sp76_16 sp77_16 11.551961
Rsn76_16 sn76_16 sn77_16 11.551961
Rsp76_17 sp76_17 sp77_17 11.551961
Rsn76_17 sn76_17 sn77_17 11.551961
Rsp76_18 sp76_18 sp77_18 11.551961
Rsn76_18 sn76_18 sn77_18 11.551961
Rsp76_19 sp76_19 sp77_19 11.551961
Rsn76_19 sn76_19 sn77_19 11.551961
Rsp76_20 sp76_20 sp77_20 11.551961
Rsn76_20 sn76_20 sn77_20 11.551961
Rsp76_21 sp76_21 sp77_21 11.551961
Rsn76_21 sn76_21 sn77_21 11.551961
Rsp76_22 sp76_22 sp77_22 11.551961
Rsn76_22 sn76_22 sn77_22 11.551961
Rsp76_23 sp76_23 sp77_23 11.551961
Rsn76_23 sn76_23 sn77_23 11.551961
Rsp76_24 sp76_24 sp77_24 11.551961
Rsn76_24 sn76_24 sn77_24 11.551961
Rsp76_25 sp76_25 sp77_25 11.551961
Rsn76_25 sn76_25 sn77_25 11.551961
Rsp76_26 sp76_26 sp77_26 11.551961
Rsn76_26 sn76_26 sn77_26 11.551961
Rsp76_27 sp76_27 sp77_27 11.551961
Rsn76_27 sn76_27 sn77_27 11.551961
Rsp76_28 sp76_28 sp77_28 11.551961
Rsn76_28 sn76_28 sn77_28 11.551961
Rsp76_29 sp76_29 sp77_29 11.551961
Rsn76_29 sn76_29 sn77_29 11.551961
Rsp76_30 sp76_30 sp77_30 11.551961
Rsn76_30 sn76_30 sn77_30 11.551961
Rsp76_31 sp76_31 sp77_31 11.551961
Rsn76_31 sn76_31 sn77_31 11.551961
Rsp76_32 sp76_32 sp77_32 11.551961
Rsn76_32 sn76_32 sn77_32 11.551961
Rsp76_33 sp76_33 sp77_33 11.551961
Rsn76_33 sn76_33 sn77_33 11.551961
Rsp76_34 sp76_34 sp77_34 11.551961
Rsn76_34 sn76_34 sn77_34 11.551961
Rsp76_35 sp76_35 sp77_35 11.551961
Rsn76_35 sn76_35 sn77_35 11.551961
Rsp76_36 sp76_36 sp77_36 11.551961
Rsn76_36 sn76_36 sn77_36 11.551961
Rsp76_37 sp76_37 sp77_37 11.551961
Rsn76_37 sn76_37 sn77_37 11.551961
Rsp76_38 sp76_38 sp77_38 11.551961
Rsn76_38 sn76_38 sn77_38 11.551961
Rsp76_39 sp76_39 sp77_39 11.551961
Rsn76_39 sn76_39 sn77_39 11.551961
Rsp76_40 sp76_40 sp77_40 11.551961
Rsn76_40 sn76_40 sn77_40 11.551961
Rsp76_41 sp76_41 sp77_41 11.551961
Rsn76_41 sn76_41 sn77_41 11.551961
Rsp76_42 sp76_42 sp77_42 11.551961
Rsn76_42 sn76_42 sn77_42 11.551961
Rsp76_43 sp76_43 sp77_43 11.551961
Rsn76_43 sn76_43 sn77_43 11.551961
Rsp76_44 sp76_44 sp77_44 11.551961
Rsn76_44 sn76_44 sn77_44 11.551961
Rsp76_45 sp76_45 sp77_45 11.551961
Rsn76_45 sn76_45 sn77_45 11.551961
Rsp76_46 sp76_46 sp77_46 11.551961
Rsn76_46 sn76_46 sn77_46 11.551961
Rsp76_47 sp76_47 sp77_47 11.551961
Rsn76_47 sn76_47 sn77_47 11.551961
Rsp76_48 sp76_48 sp77_48 11.551961
Rsn76_48 sn76_48 sn77_48 11.551961
Rsp76_49 sp76_49 sp77_49 11.551961
Rsn76_49 sn76_49 sn77_49 11.551961
Rsp76_50 sp76_50 sp77_50 11.551961
Rsn76_50 sn76_50 sn77_50 11.551961
Rsp76_51 sp76_51 sp77_51 11.551961
Rsn76_51 sn76_51 sn77_51 11.551961
Rsp76_52 sp76_52 sp77_52 11.551961
Rsn76_52 sn76_52 sn77_52 11.551961
Rsp76_53 sp76_53 sp77_53 11.551961
Rsn76_53 sn76_53 sn77_53 11.551961
Rsp76_54 sp76_54 sp77_54 11.551961
Rsn76_54 sn76_54 sn77_54 11.551961
Rsp76_55 sp76_55 sp77_55 11.551961
Rsn76_55 sn76_55 sn77_55 11.551961
Rsp76_56 sp76_56 sp77_56 11.551961
Rsn76_56 sn76_56 sn77_56 11.551961
Rsp76_57 sp76_57 sp77_57 11.551961
Rsn76_57 sn76_57 sn77_57 11.551961
Rsp76_58 sp76_58 sp77_58 11.551961
Rsn76_58 sn76_58 sn77_58 11.551961
Rsp76_59 sp76_59 sp77_59 11.551961
Rsn76_59 sn76_59 sn77_59 11.551961
Rsp76_60 sp76_60 sp77_60 11.551961
Rsn76_60 sn76_60 sn77_60 11.551961
Rsp76_61 sp76_61 sp77_61 11.551961
Rsn76_61 sn76_61 sn77_61 11.551961
Rsp76_62 sp76_62 sp77_62 11.551961
Rsn76_62 sn76_62 sn77_62 11.551961
Rsp76_63 sp76_63 sp77_63 11.551961
Rsn76_63 sn76_63 sn77_63 11.551961
Rsp76_64 sp76_64 sp77_64 11.551961
Rsn76_64 sn76_64 sn77_64 11.551961
Rsp76_65 sp76_65 sp77_65 11.551961
Rsn76_65 sn76_65 sn77_65 11.551961
Rsp76_66 sp76_66 sp77_66 11.551961
Rsn76_66 sn76_66 sn77_66 11.551961
Rsp76_67 sp76_67 sp77_67 11.551961
Rsn76_67 sn76_67 sn77_67 11.551961
Rsp76_68 sp76_68 sp77_68 11.551961
Rsn76_68 sn76_68 sn77_68 11.551961
Rsp76_69 sp76_69 sp77_69 11.551961
Rsn76_69 sn76_69 sn77_69 11.551961
Rsp76_70 sp76_70 sp77_70 11.551961
Rsn76_70 sn76_70 sn77_70 11.551961
Rsp76_71 sp76_71 sp77_71 11.551961
Rsn76_71 sn76_71 sn77_71 11.551961
Rsp76_72 sp76_72 sp77_72 11.551961
Rsn76_72 sn76_72 sn77_72 11.551961
Rsp76_73 sp76_73 sp77_73 11.551961
Rsn76_73 sn76_73 sn77_73 11.551961
Rsp76_74 sp76_74 sp77_74 11.551961
Rsn76_74 sn76_74 sn77_74 11.551961
Rsp76_75 sp76_75 sp77_75 11.551961
Rsn76_75 sn76_75 sn77_75 11.551961
Rsp76_76 sp76_76 sp77_76 11.551961
Rsn76_76 sn76_76 sn77_76 11.551961
Rsp76_77 sp76_77 sp77_77 11.551961
Rsn76_77 sn76_77 sn77_77 11.551961
Rsp76_78 sp76_78 sp77_78 11.551961
Rsn76_78 sn76_78 sn77_78 11.551961
Rsp76_79 sp76_79 sp77_79 11.551961
Rsn76_79 sn76_79 sn77_79 11.551961
Rsp76_80 sp76_80 sp77_80 11.551961
Rsn76_80 sn76_80 sn77_80 11.551961
Rsp76_81 sp76_81 sp77_81 11.551961
Rsn76_81 sn76_81 sn77_81 11.551961
Rsp76_82 sp76_82 sp77_82 11.551961
Rsn76_82 sn76_82 sn77_82 11.551961
Rsp76_83 sp76_83 sp77_83 11.551961
Rsn76_83 sn76_83 sn77_83 11.551961
Rsp76_84 sp76_84 sp77_84 11.551961
Rsn76_84 sn76_84 sn77_84 11.551961
Rsp77_1 sp77_1 sp78_1 11.551961
Rsn77_1 sn77_1 sn78_1 11.551961
Rsp77_2 sp77_2 sp78_2 11.551961
Rsn77_2 sn77_2 sn78_2 11.551961
Rsp77_3 sp77_3 sp78_3 11.551961
Rsn77_3 sn77_3 sn78_3 11.551961
Rsp77_4 sp77_4 sp78_4 11.551961
Rsn77_4 sn77_4 sn78_4 11.551961
Rsp77_5 sp77_5 sp78_5 11.551961
Rsn77_5 sn77_5 sn78_5 11.551961
Rsp77_6 sp77_6 sp78_6 11.551961
Rsn77_6 sn77_6 sn78_6 11.551961
Rsp77_7 sp77_7 sp78_7 11.551961
Rsn77_7 sn77_7 sn78_7 11.551961
Rsp77_8 sp77_8 sp78_8 11.551961
Rsn77_8 sn77_8 sn78_8 11.551961
Rsp77_9 sp77_9 sp78_9 11.551961
Rsn77_9 sn77_9 sn78_9 11.551961
Rsp77_10 sp77_10 sp78_10 11.551961
Rsn77_10 sn77_10 sn78_10 11.551961
Rsp77_11 sp77_11 sp78_11 11.551961
Rsn77_11 sn77_11 sn78_11 11.551961
Rsp77_12 sp77_12 sp78_12 11.551961
Rsn77_12 sn77_12 sn78_12 11.551961
Rsp77_13 sp77_13 sp78_13 11.551961
Rsn77_13 sn77_13 sn78_13 11.551961
Rsp77_14 sp77_14 sp78_14 11.551961
Rsn77_14 sn77_14 sn78_14 11.551961
Rsp77_15 sp77_15 sp78_15 11.551961
Rsn77_15 sn77_15 sn78_15 11.551961
Rsp77_16 sp77_16 sp78_16 11.551961
Rsn77_16 sn77_16 sn78_16 11.551961
Rsp77_17 sp77_17 sp78_17 11.551961
Rsn77_17 sn77_17 sn78_17 11.551961
Rsp77_18 sp77_18 sp78_18 11.551961
Rsn77_18 sn77_18 sn78_18 11.551961
Rsp77_19 sp77_19 sp78_19 11.551961
Rsn77_19 sn77_19 sn78_19 11.551961
Rsp77_20 sp77_20 sp78_20 11.551961
Rsn77_20 sn77_20 sn78_20 11.551961
Rsp77_21 sp77_21 sp78_21 11.551961
Rsn77_21 sn77_21 sn78_21 11.551961
Rsp77_22 sp77_22 sp78_22 11.551961
Rsn77_22 sn77_22 sn78_22 11.551961
Rsp77_23 sp77_23 sp78_23 11.551961
Rsn77_23 sn77_23 sn78_23 11.551961
Rsp77_24 sp77_24 sp78_24 11.551961
Rsn77_24 sn77_24 sn78_24 11.551961
Rsp77_25 sp77_25 sp78_25 11.551961
Rsn77_25 sn77_25 sn78_25 11.551961
Rsp77_26 sp77_26 sp78_26 11.551961
Rsn77_26 sn77_26 sn78_26 11.551961
Rsp77_27 sp77_27 sp78_27 11.551961
Rsn77_27 sn77_27 sn78_27 11.551961
Rsp77_28 sp77_28 sp78_28 11.551961
Rsn77_28 sn77_28 sn78_28 11.551961
Rsp77_29 sp77_29 sp78_29 11.551961
Rsn77_29 sn77_29 sn78_29 11.551961
Rsp77_30 sp77_30 sp78_30 11.551961
Rsn77_30 sn77_30 sn78_30 11.551961
Rsp77_31 sp77_31 sp78_31 11.551961
Rsn77_31 sn77_31 sn78_31 11.551961
Rsp77_32 sp77_32 sp78_32 11.551961
Rsn77_32 sn77_32 sn78_32 11.551961
Rsp77_33 sp77_33 sp78_33 11.551961
Rsn77_33 sn77_33 sn78_33 11.551961
Rsp77_34 sp77_34 sp78_34 11.551961
Rsn77_34 sn77_34 sn78_34 11.551961
Rsp77_35 sp77_35 sp78_35 11.551961
Rsn77_35 sn77_35 sn78_35 11.551961
Rsp77_36 sp77_36 sp78_36 11.551961
Rsn77_36 sn77_36 sn78_36 11.551961
Rsp77_37 sp77_37 sp78_37 11.551961
Rsn77_37 sn77_37 sn78_37 11.551961
Rsp77_38 sp77_38 sp78_38 11.551961
Rsn77_38 sn77_38 sn78_38 11.551961
Rsp77_39 sp77_39 sp78_39 11.551961
Rsn77_39 sn77_39 sn78_39 11.551961
Rsp77_40 sp77_40 sp78_40 11.551961
Rsn77_40 sn77_40 sn78_40 11.551961
Rsp77_41 sp77_41 sp78_41 11.551961
Rsn77_41 sn77_41 sn78_41 11.551961
Rsp77_42 sp77_42 sp78_42 11.551961
Rsn77_42 sn77_42 sn78_42 11.551961
Rsp77_43 sp77_43 sp78_43 11.551961
Rsn77_43 sn77_43 sn78_43 11.551961
Rsp77_44 sp77_44 sp78_44 11.551961
Rsn77_44 sn77_44 sn78_44 11.551961
Rsp77_45 sp77_45 sp78_45 11.551961
Rsn77_45 sn77_45 sn78_45 11.551961
Rsp77_46 sp77_46 sp78_46 11.551961
Rsn77_46 sn77_46 sn78_46 11.551961
Rsp77_47 sp77_47 sp78_47 11.551961
Rsn77_47 sn77_47 sn78_47 11.551961
Rsp77_48 sp77_48 sp78_48 11.551961
Rsn77_48 sn77_48 sn78_48 11.551961
Rsp77_49 sp77_49 sp78_49 11.551961
Rsn77_49 sn77_49 sn78_49 11.551961
Rsp77_50 sp77_50 sp78_50 11.551961
Rsn77_50 sn77_50 sn78_50 11.551961
Rsp77_51 sp77_51 sp78_51 11.551961
Rsn77_51 sn77_51 sn78_51 11.551961
Rsp77_52 sp77_52 sp78_52 11.551961
Rsn77_52 sn77_52 sn78_52 11.551961
Rsp77_53 sp77_53 sp78_53 11.551961
Rsn77_53 sn77_53 sn78_53 11.551961
Rsp77_54 sp77_54 sp78_54 11.551961
Rsn77_54 sn77_54 sn78_54 11.551961
Rsp77_55 sp77_55 sp78_55 11.551961
Rsn77_55 sn77_55 sn78_55 11.551961
Rsp77_56 sp77_56 sp78_56 11.551961
Rsn77_56 sn77_56 sn78_56 11.551961
Rsp77_57 sp77_57 sp78_57 11.551961
Rsn77_57 sn77_57 sn78_57 11.551961
Rsp77_58 sp77_58 sp78_58 11.551961
Rsn77_58 sn77_58 sn78_58 11.551961
Rsp77_59 sp77_59 sp78_59 11.551961
Rsn77_59 sn77_59 sn78_59 11.551961
Rsp77_60 sp77_60 sp78_60 11.551961
Rsn77_60 sn77_60 sn78_60 11.551961
Rsp77_61 sp77_61 sp78_61 11.551961
Rsn77_61 sn77_61 sn78_61 11.551961
Rsp77_62 sp77_62 sp78_62 11.551961
Rsn77_62 sn77_62 sn78_62 11.551961
Rsp77_63 sp77_63 sp78_63 11.551961
Rsn77_63 sn77_63 sn78_63 11.551961
Rsp77_64 sp77_64 sp78_64 11.551961
Rsn77_64 sn77_64 sn78_64 11.551961
Rsp77_65 sp77_65 sp78_65 11.551961
Rsn77_65 sn77_65 sn78_65 11.551961
Rsp77_66 sp77_66 sp78_66 11.551961
Rsn77_66 sn77_66 sn78_66 11.551961
Rsp77_67 sp77_67 sp78_67 11.551961
Rsn77_67 sn77_67 sn78_67 11.551961
Rsp77_68 sp77_68 sp78_68 11.551961
Rsn77_68 sn77_68 sn78_68 11.551961
Rsp77_69 sp77_69 sp78_69 11.551961
Rsn77_69 sn77_69 sn78_69 11.551961
Rsp77_70 sp77_70 sp78_70 11.551961
Rsn77_70 sn77_70 sn78_70 11.551961
Rsp77_71 sp77_71 sp78_71 11.551961
Rsn77_71 sn77_71 sn78_71 11.551961
Rsp77_72 sp77_72 sp78_72 11.551961
Rsn77_72 sn77_72 sn78_72 11.551961
Rsp77_73 sp77_73 sp78_73 11.551961
Rsn77_73 sn77_73 sn78_73 11.551961
Rsp77_74 sp77_74 sp78_74 11.551961
Rsn77_74 sn77_74 sn78_74 11.551961
Rsp77_75 sp77_75 sp78_75 11.551961
Rsn77_75 sn77_75 sn78_75 11.551961
Rsp77_76 sp77_76 sp78_76 11.551961
Rsn77_76 sn77_76 sn78_76 11.551961
Rsp77_77 sp77_77 sp78_77 11.551961
Rsn77_77 sn77_77 sn78_77 11.551961
Rsp77_78 sp77_78 sp78_78 11.551961
Rsn77_78 sn77_78 sn78_78 11.551961
Rsp77_79 sp77_79 sp78_79 11.551961
Rsn77_79 sn77_79 sn78_79 11.551961
Rsp77_80 sp77_80 sp78_80 11.551961
Rsn77_80 sn77_80 sn78_80 11.551961
Rsp77_81 sp77_81 sp78_81 11.551961
Rsn77_81 sn77_81 sn78_81 11.551961
Rsp77_82 sp77_82 sp78_82 11.551961
Rsn77_82 sn77_82 sn78_82 11.551961
Rsp77_83 sp77_83 sp78_83 11.551961
Rsn77_83 sn77_83 sn78_83 11.551961
Rsp77_84 sp77_84 sp78_84 11.551961
Rsn77_84 sn77_84 sn78_84 11.551961
Rsp78_1 sp78_1 sp79_1 11.551961
Rsn78_1 sn78_1 sn79_1 11.551961
Rsp78_2 sp78_2 sp79_2 11.551961
Rsn78_2 sn78_2 sn79_2 11.551961
Rsp78_3 sp78_3 sp79_3 11.551961
Rsn78_3 sn78_3 sn79_3 11.551961
Rsp78_4 sp78_4 sp79_4 11.551961
Rsn78_4 sn78_4 sn79_4 11.551961
Rsp78_5 sp78_5 sp79_5 11.551961
Rsn78_5 sn78_5 sn79_5 11.551961
Rsp78_6 sp78_6 sp79_6 11.551961
Rsn78_6 sn78_6 sn79_6 11.551961
Rsp78_7 sp78_7 sp79_7 11.551961
Rsn78_7 sn78_7 sn79_7 11.551961
Rsp78_8 sp78_8 sp79_8 11.551961
Rsn78_8 sn78_8 sn79_8 11.551961
Rsp78_9 sp78_9 sp79_9 11.551961
Rsn78_9 sn78_9 sn79_9 11.551961
Rsp78_10 sp78_10 sp79_10 11.551961
Rsn78_10 sn78_10 sn79_10 11.551961
Rsp78_11 sp78_11 sp79_11 11.551961
Rsn78_11 sn78_11 sn79_11 11.551961
Rsp78_12 sp78_12 sp79_12 11.551961
Rsn78_12 sn78_12 sn79_12 11.551961
Rsp78_13 sp78_13 sp79_13 11.551961
Rsn78_13 sn78_13 sn79_13 11.551961
Rsp78_14 sp78_14 sp79_14 11.551961
Rsn78_14 sn78_14 sn79_14 11.551961
Rsp78_15 sp78_15 sp79_15 11.551961
Rsn78_15 sn78_15 sn79_15 11.551961
Rsp78_16 sp78_16 sp79_16 11.551961
Rsn78_16 sn78_16 sn79_16 11.551961
Rsp78_17 sp78_17 sp79_17 11.551961
Rsn78_17 sn78_17 sn79_17 11.551961
Rsp78_18 sp78_18 sp79_18 11.551961
Rsn78_18 sn78_18 sn79_18 11.551961
Rsp78_19 sp78_19 sp79_19 11.551961
Rsn78_19 sn78_19 sn79_19 11.551961
Rsp78_20 sp78_20 sp79_20 11.551961
Rsn78_20 sn78_20 sn79_20 11.551961
Rsp78_21 sp78_21 sp79_21 11.551961
Rsn78_21 sn78_21 sn79_21 11.551961
Rsp78_22 sp78_22 sp79_22 11.551961
Rsn78_22 sn78_22 sn79_22 11.551961
Rsp78_23 sp78_23 sp79_23 11.551961
Rsn78_23 sn78_23 sn79_23 11.551961
Rsp78_24 sp78_24 sp79_24 11.551961
Rsn78_24 sn78_24 sn79_24 11.551961
Rsp78_25 sp78_25 sp79_25 11.551961
Rsn78_25 sn78_25 sn79_25 11.551961
Rsp78_26 sp78_26 sp79_26 11.551961
Rsn78_26 sn78_26 sn79_26 11.551961
Rsp78_27 sp78_27 sp79_27 11.551961
Rsn78_27 sn78_27 sn79_27 11.551961
Rsp78_28 sp78_28 sp79_28 11.551961
Rsn78_28 sn78_28 sn79_28 11.551961
Rsp78_29 sp78_29 sp79_29 11.551961
Rsn78_29 sn78_29 sn79_29 11.551961
Rsp78_30 sp78_30 sp79_30 11.551961
Rsn78_30 sn78_30 sn79_30 11.551961
Rsp78_31 sp78_31 sp79_31 11.551961
Rsn78_31 sn78_31 sn79_31 11.551961
Rsp78_32 sp78_32 sp79_32 11.551961
Rsn78_32 sn78_32 sn79_32 11.551961
Rsp78_33 sp78_33 sp79_33 11.551961
Rsn78_33 sn78_33 sn79_33 11.551961
Rsp78_34 sp78_34 sp79_34 11.551961
Rsn78_34 sn78_34 sn79_34 11.551961
Rsp78_35 sp78_35 sp79_35 11.551961
Rsn78_35 sn78_35 sn79_35 11.551961
Rsp78_36 sp78_36 sp79_36 11.551961
Rsn78_36 sn78_36 sn79_36 11.551961
Rsp78_37 sp78_37 sp79_37 11.551961
Rsn78_37 sn78_37 sn79_37 11.551961
Rsp78_38 sp78_38 sp79_38 11.551961
Rsn78_38 sn78_38 sn79_38 11.551961
Rsp78_39 sp78_39 sp79_39 11.551961
Rsn78_39 sn78_39 sn79_39 11.551961
Rsp78_40 sp78_40 sp79_40 11.551961
Rsn78_40 sn78_40 sn79_40 11.551961
Rsp78_41 sp78_41 sp79_41 11.551961
Rsn78_41 sn78_41 sn79_41 11.551961
Rsp78_42 sp78_42 sp79_42 11.551961
Rsn78_42 sn78_42 sn79_42 11.551961
Rsp78_43 sp78_43 sp79_43 11.551961
Rsn78_43 sn78_43 sn79_43 11.551961
Rsp78_44 sp78_44 sp79_44 11.551961
Rsn78_44 sn78_44 sn79_44 11.551961
Rsp78_45 sp78_45 sp79_45 11.551961
Rsn78_45 sn78_45 sn79_45 11.551961
Rsp78_46 sp78_46 sp79_46 11.551961
Rsn78_46 sn78_46 sn79_46 11.551961
Rsp78_47 sp78_47 sp79_47 11.551961
Rsn78_47 sn78_47 sn79_47 11.551961
Rsp78_48 sp78_48 sp79_48 11.551961
Rsn78_48 sn78_48 sn79_48 11.551961
Rsp78_49 sp78_49 sp79_49 11.551961
Rsn78_49 sn78_49 sn79_49 11.551961
Rsp78_50 sp78_50 sp79_50 11.551961
Rsn78_50 sn78_50 sn79_50 11.551961
Rsp78_51 sp78_51 sp79_51 11.551961
Rsn78_51 sn78_51 sn79_51 11.551961
Rsp78_52 sp78_52 sp79_52 11.551961
Rsn78_52 sn78_52 sn79_52 11.551961
Rsp78_53 sp78_53 sp79_53 11.551961
Rsn78_53 sn78_53 sn79_53 11.551961
Rsp78_54 sp78_54 sp79_54 11.551961
Rsn78_54 sn78_54 sn79_54 11.551961
Rsp78_55 sp78_55 sp79_55 11.551961
Rsn78_55 sn78_55 sn79_55 11.551961
Rsp78_56 sp78_56 sp79_56 11.551961
Rsn78_56 sn78_56 sn79_56 11.551961
Rsp78_57 sp78_57 sp79_57 11.551961
Rsn78_57 sn78_57 sn79_57 11.551961
Rsp78_58 sp78_58 sp79_58 11.551961
Rsn78_58 sn78_58 sn79_58 11.551961
Rsp78_59 sp78_59 sp79_59 11.551961
Rsn78_59 sn78_59 sn79_59 11.551961
Rsp78_60 sp78_60 sp79_60 11.551961
Rsn78_60 sn78_60 sn79_60 11.551961
Rsp78_61 sp78_61 sp79_61 11.551961
Rsn78_61 sn78_61 sn79_61 11.551961
Rsp78_62 sp78_62 sp79_62 11.551961
Rsn78_62 sn78_62 sn79_62 11.551961
Rsp78_63 sp78_63 sp79_63 11.551961
Rsn78_63 sn78_63 sn79_63 11.551961
Rsp78_64 sp78_64 sp79_64 11.551961
Rsn78_64 sn78_64 sn79_64 11.551961
Rsp78_65 sp78_65 sp79_65 11.551961
Rsn78_65 sn78_65 sn79_65 11.551961
Rsp78_66 sp78_66 sp79_66 11.551961
Rsn78_66 sn78_66 sn79_66 11.551961
Rsp78_67 sp78_67 sp79_67 11.551961
Rsn78_67 sn78_67 sn79_67 11.551961
Rsp78_68 sp78_68 sp79_68 11.551961
Rsn78_68 sn78_68 sn79_68 11.551961
Rsp78_69 sp78_69 sp79_69 11.551961
Rsn78_69 sn78_69 sn79_69 11.551961
Rsp78_70 sp78_70 sp79_70 11.551961
Rsn78_70 sn78_70 sn79_70 11.551961
Rsp78_71 sp78_71 sp79_71 11.551961
Rsn78_71 sn78_71 sn79_71 11.551961
Rsp78_72 sp78_72 sp79_72 11.551961
Rsn78_72 sn78_72 sn79_72 11.551961
Rsp78_73 sp78_73 sp79_73 11.551961
Rsn78_73 sn78_73 sn79_73 11.551961
Rsp78_74 sp78_74 sp79_74 11.551961
Rsn78_74 sn78_74 sn79_74 11.551961
Rsp78_75 sp78_75 sp79_75 11.551961
Rsn78_75 sn78_75 sn79_75 11.551961
Rsp78_76 sp78_76 sp79_76 11.551961
Rsn78_76 sn78_76 sn79_76 11.551961
Rsp78_77 sp78_77 sp79_77 11.551961
Rsn78_77 sn78_77 sn79_77 11.551961
Rsp78_78 sp78_78 sp79_78 11.551961
Rsn78_78 sn78_78 sn79_78 11.551961
Rsp78_79 sp78_79 sp79_79 11.551961
Rsn78_79 sn78_79 sn79_79 11.551961
Rsp78_80 sp78_80 sp79_80 11.551961
Rsn78_80 sn78_80 sn79_80 11.551961
Rsp78_81 sp78_81 sp79_81 11.551961
Rsn78_81 sn78_81 sn79_81 11.551961
Rsp78_82 sp78_82 sp79_82 11.551961
Rsn78_82 sn78_82 sn79_82 11.551961
Rsp78_83 sp78_83 sp79_83 11.551961
Rsn78_83 sn78_83 sn79_83 11.551961
Rsp78_84 sp78_84 sp79_84 11.551961
Rsn78_84 sn78_84 sn79_84 11.551961
Rsp79_1 sp79_1 sp80_1 11.551961
Rsn79_1 sn79_1 sn80_1 11.551961
Rsp79_2 sp79_2 sp80_2 11.551961
Rsn79_2 sn79_2 sn80_2 11.551961
Rsp79_3 sp79_3 sp80_3 11.551961
Rsn79_3 sn79_3 sn80_3 11.551961
Rsp79_4 sp79_4 sp80_4 11.551961
Rsn79_4 sn79_4 sn80_4 11.551961
Rsp79_5 sp79_5 sp80_5 11.551961
Rsn79_5 sn79_5 sn80_5 11.551961
Rsp79_6 sp79_6 sp80_6 11.551961
Rsn79_6 sn79_6 sn80_6 11.551961
Rsp79_7 sp79_7 sp80_7 11.551961
Rsn79_7 sn79_7 sn80_7 11.551961
Rsp79_8 sp79_8 sp80_8 11.551961
Rsn79_8 sn79_8 sn80_8 11.551961
Rsp79_9 sp79_9 sp80_9 11.551961
Rsn79_9 sn79_9 sn80_9 11.551961
Rsp79_10 sp79_10 sp80_10 11.551961
Rsn79_10 sn79_10 sn80_10 11.551961
Rsp79_11 sp79_11 sp80_11 11.551961
Rsn79_11 sn79_11 sn80_11 11.551961
Rsp79_12 sp79_12 sp80_12 11.551961
Rsn79_12 sn79_12 sn80_12 11.551961
Rsp79_13 sp79_13 sp80_13 11.551961
Rsn79_13 sn79_13 sn80_13 11.551961
Rsp79_14 sp79_14 sp80_14 11.551961
Rsn79_14 sn79_14 sn80_14 11.551961
Rsp79_15 sp79_15 sp80_15 11.551961
Rsn79_15 sn79_15 sn80_15 11.551961
Rsp79_16 sp79_16 sp80_16 11.551961
Rsn79_16 sn79_16 sn80_16 11.551961
Rsp79_17 sp79_17 sp80_17 11.551961
Rsn79_17 sn79_17 sn80_17 11.551961
Rsp79_18 sp79_18 sp80_18 11.551961
Rsn79_18 sn79_18 sn80_18 11.551961
Rsp79_19 sp79_19 sp80_19 11.551961
Rsn79_19 sn79_19 sn80_19 11.551961
Rsp79_20 sp79_20 sp80_20 11.551961
Rsn79_20 sn79_20 sn80_20 11.551961
Rsp79_21 sp79_21 sp80_21 11.551961
Rsn79_21 sn79_21 sn80_21 11.551961
Rsp79_22 sp79_22 sp80_22 11.551961
Rsn79_22 sn79_22 sn80_22 11.551961
Rsp79_23 sp79_23 sp80_23 11.551961
Rsn79_23 sn79_23 sn80_23 11.551961
Rsp79_24 sp79_24 sp80_24 11.551961
Rsn79_24 sn79_24 sn80_24 11.551961
Rsp79_25 sp79_25 sp80_25 11.551961
Rsn79_25 sn79_25 sn80_25 11.551961
Rsp79_26 sp79_26 sp80_26 11.551961
Rsn79_26 sn79_26 sn80_26 11.551961
Rsp79_27 sp79_27 sp80_27 11.551961
Rsn79_27 sn79_27 sn80_27 11.551961
Rsp79_28 sp79_28 sp80_28 11.551961
Rsn79_28 sn79_28 sn80_28 11.551961
Rsp79_29 sp79_29 sp80_29 11.551961
Rsn79_29 sn79_29 sn80_29 11.551961
Rsp79_30 sp79_30 sp80_30 11.551961
Rsn79_30 sn79_30 sn80_30 11.551961
Rsp79_31 sp79_31 sp80_31 11.551961
Rsn79_31 sn79_31 sn80_31 11.551961
Rsp79_32 sp79_32 sp80_32 11.551961
Rsn79_32 sn79_32 sn80_32 11.551961
Rsp79_33 sp79_33 sp80_33 11.551961
Rsn79_33 sn79_33 sn80_33 11.551961
Rsp79_34 sp79_34 sp80_34 11.551961
Rsn79_34 sn79_34 sn80_34 11.551961
Rsp79_35 sp79_35 sp80_35 11.551961
Rsn79_35 sn79_35 sn80_35 11.551961
Rsp79_36 sp79_36 sp80_36 11.551961
Rsn79_36 sn79_36 sn80_36 11.551961
Rsp79_37 sp79_37 sp80_37 11.551961
Rsn79_37 sn79_37 sn80_37 11.551961
Rsp79_38 sp79_38 sp80_38 11.551961
Rsn79_38 sn79_38 sn80_38 11.551961
Rsp79_39 sp79_39 sp80_39 11.551961
Rsn79_39 sn79_39 sn80_39 11.551961
Rsp79_40 sp79_40 sp80_40 11.551961
Rsn79_40 sn79_40 sn80_40 11.551961
Rsp79_41 sp79_41 sp80_41 11.551961
Rsn79_41 sn79_41 sn80_41 11.551961
Rsp79_42 sp79_42 sp80_42 11.551961
Rsn79_42 sn79_42 sn80_42 11.551961
Rsp79_43 sp79_43 sp80_43 11.551961
Rsn79_43 sn79_43 sn80_43 11.551961
Rsp79_44 sp79_44 sp80_44 11.551961
Rsn79_44 sn79_44 sn80_44 11.551961
Rsp79_45 sp79_45 sp80_45 11.551961
Rsn79_45 sn79_45 sn80_45 11.551961
Rsp79_46 sp79_46 sp80_46 11.551961
Rsn79_46 sn79_46 sn80_46 11.551961
Rsp79_47 sp79_47 sp80_47 11.551961
Rsn79_47 sn79_47 sn80_47 11.551961
Rsp79_48 sp79_48 sp80_48 11.551961
Rsn79_48 sn79_48 sn80_48 11.551961
Rsp79_49 sp79_49 sp80_49 11.551961
Rsn79_49 sn79_49 sn80_49 11.551961
Rsp79_50 sp79_50 sp80_50 11.551961
Rsn79_50 sn79_50 sn80_50 11.551961
Rsp79_51 sp79_51 sp80_51 11.551961
Rsn79_51 sn79_51 sn80_51 11.551961
Rsp79_52 sp79_52 sp80_52 11.551961
Rsn79_52 sn79_52 sn80_52 11.551961
Rsp79_53 sp79_53 sp80_53 11.551961
Rsn79_53 sn79_53 sn80_53 11.551961
Rsp79_54 sp79_54 sp80_54 11.551961
Rsn79_54 sn79_54 sn80_54 11.551961
Rsp79_55 sp79_55 sp80_55 11.551961
Rsn79_55 sn79_55 sn80_55 11.551961
Rsp79_56 sp79_56 sp80_56 11.551961
Rsn79_56 sn79_56 sn80_56 11.551961
Rsp79_57 sp79_57 sp80_57 11.551961
Rsn79_57 sn79_57 sn80_57 11.551961
Rsp79_58 sp79_58 sp80_58 11.551961
Rsn79_58 sn79_58 sn80_58 11.551961
Rsp79_59 sp79_59 sp80_59 11.551961
Rsn79_59 sn79_59 sn80_59 11.551961
Rsp79_60 sp79_60 sp80_60 11.551961
Rsn79_60 sn79_60 sn80_60 11.551961
Rsp79_61 sp79_61 sp80_61 11.551961
Rsn79_61 sn79_61 sn80_61 11.551961
Rsp79_62 sp79_62 sp80_62 11.551961
Rsn79_62 sn79_62 sn80_62 11.551961
Rsp79_63 sp79_63 sp80_63 11.551961
Rsn79_63 sn79_63 sn80_63 11.551961
Rsp79_64 sp79_64 sp80_64 11.551961
Rsn79_64 sn79_64 sn80_64 11.551961
Rsp79_65 sp79_65 sp80_65 11.551961
Rsn79_65 sn79_65 sn80_65 11.551961
Rsp79_66 sp79_66 sp80_66 11.551961
Rsn79_66 sn79_66 sn80_66 11.551961
Rsp79_67 sp79_67 sp80_67 11.551961
Rsn79_67 sn79_67 sn80_67 11.551961
Rsp79_68 sp79_68 sp80_68 11.551961
Rsn79_68 sn79_68 sn80_68 11.551961
Rsp79_69 sp79_69 sp80_69 11.551961
Rsn79_69 sn79_69 sn80_69 11.551961
Rsp79_70 sp79_70 sp80_70 11.551961
Rsn79_70 sn79_70 sn80_70 11.551961
Rsp79_71 sp79_71 sp80_71 11.551961
Rsn79_71 sn79_71 sn80_71 11.551961
Rsp79_72 sp79_72 sp80_72 11.551961
Rsn79_72 sn79_72 sn80_72 11.551961
Rsp79_73 sp79_73 sp80_73 11.551961
Rsn79_73 sn79_73 sn80_73 11.551961
Rsp79_74 sp79_74 sp80_74 11.551961
Rsn79_74 sn79_74 sn80_74 11.551961
Rsp79_75 sp79_75 sp80_75 11.551961
Rsn79_75 sn79_75 sn80_75 11.551961
Rsp79_76 sp79_76 sp80_76 11.551961
Rsn79_76 sn79_76 sn80_76 11.551961
Rsp79_77 sp79_77 sp80_77 11.551961
Rsn79_77 sn79_77 sn80_77 11.551961
Rsp79_78 sp79_78 sp80_78 11.551961
Rsn79_78 sn79_78 sn80_78 11.551961
Rsp79_79 sp79_79 sp80_79 11.551961
Rsn79_79 sn79_79 sn80_79 11.551961
Rsp79_80 sp79_80 sp80_80 11.551961
Rsn79_80 sn79_80 sn80_80 11.551961
Rsp79_81 sp79_81 sp80_81 11.551961
Rsn79_81 sn79_81 sn80_81 11.551961
Rsp79_82 sp79_82 sp80_82 11.551961
Rsn79_82 sn79_82 sn80_82 11.551961
Rsp79_83 sp79_83 sp80_83 11.551961
Rsn79_83 sn79_83 sn80_83 11.551961
Rsp79_84 sp79_84 sp80_84 11.551961
Rsn79_84 sn79_84 sn80_84 11.551961
Rsp80_1 sp80_1 sp81_1 11.551961
Rsn80_1 sn80_1 sn81_1 11.551961
Rsp80_2 sp80_2 sp81_2 11.551961
Rsn80_2 sn80_2 sn81_2 11.551961
Rsp80_3 sp80_3 sp81_3 11.551961
Rsn80_3 sn80_3 sn81_3 11.551961
Rsp80_4 sp80_4 sp81_4 11.551961
Rsn80_4 sn80_4 sn81_4 11.551961
Rsp80_5 sp80_5 sp81_5 11.551961
Rsn80_5 sn80_5 sn81_5 11.551961
Rsp80_6 sp80_6 sp81_6 11.551961
Rsn80_6 sn80_6 sn81_6 11.551961
Rsp80_7 sp80_7 sp81_7 11.551961
Rsn80_7 sn80_7 sn81_7 11.551961
Rsp80_8 sp80_8 sp81_8 11.551961
Rsn80_8 sn80_8 sn81_8 11.551961
Rsp80_9 sp80_9 sp81_9 11.551961
Rsn80_9 sn80_9 sn81_9 11.551961
Rsp80_10 sp80_10 sp81_10 11.551961
Rsn80_10 sn80_10 sn81_10 11.551961
Rsp80_11 sp80_11 sp81_11 11.551961
Rsn80_11 sn80_11 sn81_11 11.551961
Rsp80_12 sp80_12 sp81_12 11.551961
Rsn80_12 sn80_12 sn81_12 11.551961
Rsp80_13 sp80_13 sp81_13 11.551961
Rsn80_13 sn80_13 sn81_13 11.551961
Rsp80_14 sp80_14 sp81_14 11.551961
Rsn80_14 sn80_14 sn81_14 11.551961
Rsp80_15 sp80_15 sp81_15 11.551961
Rsn80_15 sn80_15 sn81_15 11.551961
Rsp80_16 sp80_16 sp81_16 11.551961
Rsn80_16 sn80_16 sn81_16 11.551961
Rsp80_17 sp80_17 sp81_17 11.551961
Rsn80_17 sn80_17 sn81_17 11.551961
Rsp80_18 sp80_18 sp81_18 11.551961
Rsn80_18 sn80_18 sn81_18 11.551961
Rsp80_19 sp80_19 sp81_19 11.551961
Rsn80_19 sn80_19 sn81_19 11.551961
Rsp80_20 sp80_20 sp81_20 11.551961
Rsn80_20 sn80_20 sn81_20 11.551961
Rsp80_21 sp80_21 sp81_21 11.551961
Rsn80_21 sn80_21 sn81_21 11.551961
Rsp80_22 sp80_22 sp81_22 11.551961
Rsn80_22 sn80_22 sn81_22 11.551961
Rsp80_23 sp80_23 sp81_23 11.551961
Rsn80_23 sn80_23 sn81_23 11.551961
Rsp80_24 sp80_24 sp81_24 11.551961
Rsn80_24 sn80_24 sn81_24 11.551961
Rsp80_25 sp80_25 sp81_25 11.551961
Rsn80_25 sn80_25 sn81_25 11.551961
Rsp80_26 sp80_26 sp81_26 11.551961
Rsn80_26 sn80_26 sn81_26 11.551961
Rsp80_27 sp80_27 sp81_27 11.551961
Rsn80_27 sn80_27 sn81_27 11.551961
Rsp80_28 sp80_28 sp81_28 11.551961
Rsn80_28 sn80_28 sn81_28 11.551961
Rsp80_29 sp80_29 sp81_29 11.551961
Rsn80_29 sn80_29 sn81_29 11.551961
Rsp80_30 sp80_30 sp81_30 11.551961
Rsn80_30 sn80_30 sn81_30 11.551961
Rsp80_31 sp80_31 sp81_31 11.551961
Rsn80_31 sn80_31 sn81_31 11.551961
Rsp80_32 sp80_32 sp81_32 11.551961
Rsn80_32 sn80_32 sn81_32 11.551961
Rsp80_33 sp80_33 sp81_33 11.551961
Rsn80_33 sn80_33 sn81_33 11.551961
Rsp80_34 sp80_34 sp81_34 11.551961
Rsn80_34 sn80_34 sn81_34 11.551961
Rsp80_35 sp80_35 sp81_35 11.551961
Rsn80_35 sn80_35 sn81_35 11.551961
Rsp80_36 sp80_36 sp81_36 11.551961
Rsn80_36 sn80_36 sn81_36 11.551961
Rsp80_37 sp80_37 sp81_37 11.551961
Rsn80_37 sn80_37 sn81_37 11.551961
Rsp80_38 sp80_38 sp81_38 11.551961
Rsn80_38 sn80_38 sn81_38 11.551961
Rsp80_39 sp80_39 sp81_39 11.551961
Rsn80_39 sn80_39 sn81_39 11.551961
Rsp80_40 sp80_40 sp81_40 11.551961
Rsn80_40 sn80_40 sn81_40 11.551961
Rsp80_41 sp80_41 sp81_41 11.551961
Rsn80_41 sn80_41 sn81_41 11.551961
Rsp80_42 sp80_42 sp81_42 11.551961
Rsn80_42 sn80_42 sn81_42 11.551961
Rsp80_43 sp80_43 sp81_43 11.551961
Rsn80_43 sn80_43 sn81_43 11.551961
Rsp80_44 sp80_44 sp81_44 11.551961
Rsn80_44 sn80_44 sn81_44 11.551961
Rsp80_45 sp80_45 sp81_45 11.551961
Rsn80_45 sn80_45 sn81_45 11.551961
Rsp80_46 sp80_46 sp81_46 11.551961
Rsn80_46 sn80_46 sn81_46 11.551961
Rsp80_47 sp80_47 sp81_47 11.551961
Rsn80_47 sn80_47 sn81_47 11.551961
Rsp80_48 sp80_48 sp81_48 11.551961
Rsn80_48 sn80_48 sn81_48 11.551961
Rsp80_49 sp80_49 sp81_49 11.551961
Rsn80_49 sn80_49 sn81_49 11.551961
Rsp80_50 sp80_50 sp81_50 11.551961
Rsn80_50 sn80_50 sn81_50 11.551961
Rsp80_51 sp80_51 sp81_51 11.551961
Rsn80_51 sn80_51 sn81_51 11.551961
Rsp80_52 sp80_52 sp81_52 11.551961
Rsn80_52 sn80_52 sn81_52 11.551961
Rsp80_53 sp80_53 sp81_53 11.551961
Rsn80_53 sn80_53 sn81_53 11.551961
Rsp80_54 sp80_54 sp81_54 11.551961
Rsn80_54 sn80_54 sn81_54 11.551961
Rsp80_55 sp80_55 sp81_55 11.551961
Rsn80_55 sn80_55 sn81_55 11.551961
Rsp80_56 sp80_56 sp81_56 11.551961
Rsn80_56 sn80_56 sn81_56 11.551961
Rsp80_57 sp80_57 sp81_57 11.551961
Rsn80_57 sn80_57 sn81_57 11.551961
Rsp80_58 sp80_58 sp81_58 11.551961
Rsn80_58 sn80_58 sn81_58 11.551961
Rsp80_59 sp80_59 sp81_59 11.551961
Rsn80_59 sn80_59 sn81_59 11.551961
Rsp80_60 sp80_60 sp81_60 11.551961
Rsn80_60 sn80_60 sn81_60 11.551961
Rsp80_61 sp80_61 sp81_61 11.551961
Rsn80_61 sn80_61 sn81_61 11.551961
Rsp80_62 sp80_62 sp81_62 11.551961
Rsn80_62 sn80_62 sn81_62 11.551961
Rsp80_63 sp80_63 sp81_63 11.551961
Rsn80_63 sn80_63 sn81_63 11.551961
Rsp80_64 sp80_64 sp81_64 11.551961
Rsn80_64 sn80_64 sn81_64 11.551961
Rsp80_65 sp80_65 sp81_65 11.551961
Rsn80_65 sn80_65 sn81_65 11.551961
Rsp80_66 sp80_66 sp81_66 11.551961
Rsn80_66 sn80_66 sn81_66 11.551961
Rsp80_67 sp80_67 sp81_67 11.551961
Rsn80_67 sn80_67 sn81_67 11.551961
Rsp80_68 sp80_68 sp81_68 11.551961
Rsn80_68 sn80_68 sn81_68 11.551961
Rsp80_69 sp80_69 sp81_69 11.551961
Rsn80_69 sn80_69 sn81_69 11.551961
Rsp80_70 sp80_70 sp81_70 11.551961
Rsn80_70 sn80_70 sn81_70 11.551961
Rsp80_71 sp80_71 sp81_71 11.551961
Rsn80_71 sn80_71 sn81_71 11.551961
Rsp80_72 sp80_72 sp81_72 11.551961
Rsn80_72 sn80_72 sn81_72 11.551961
Rsp80_73 sp80_73 sp81_73 11.551961
Rsn80_73 sn80_73 sn81_73 11.551961
Rsp80_74 sp80_74 sp81_74 11.551961
Rsn80_74 sn80_74 sn81_74 11.551961
Rsp80_75 sp80_75 sp81_75 11.551961
Rsn80_75 sn80_75 sn81_75 11.551961
Rsp80_76 sp80_76 sp81_76 11.551961
Rsn80_76 sn80_76 sn81_76 11.551961
Rsp80_77 sp80_77 sp81_77 11.551961
Rsn80_77 sn80_77 sn81_77 11.551961
Rsp80_78 sp80_78 sp81_78 11.551961
Rsn80_78 sn80_78 sn81_78 11.551961
Rsp80_79 sp80_79 sp81_79 11.551961
Rsn80_79 sn80_79 sn81_79 11.551961
Rsp80_80 sp80_80 sp81_80 11.551961
Rsn80_80 sn80_80 sn81_80 11.551961
Rsp80_81 sp80_81 sp81_81 11.551961
Rsn80_81 sn80_81 sn81_81 11.551961
Rsp80_82 sp80_82 sp81_82 11.551961
Rsn80_82 sn80_82 sn81_82 11.551961
Rsp80_83 sp80_83 sp81_83 11.551961
Rsn80_83 sn80_83 sn81_83 11.551961
Rsp80_84 sp80_84 sp81_84 11.551961
Rsn80_84 sn80_84 sn81_84 11.551961
Rsp81_1 sp81_1 sp82_1 11.551961
Rsn81_1 sn81_1 sn82_1 11.551961
Rsp81_2 sp81_2 sp82_2 11.551961
Rsn81_2 sn81_2 sn82_2 11.551961
Rsp81_3 sp81_3 sp82_3 11.551961
Rsn81_3 sn81_3 sn82_3 11.551961
Rsp81_4 sp81_4 sp82_4 11.551961
Rsn81_4 sn81_4 sn82_4 11.551961
Rsp81_5 sp81_5 sp82_5 11.551961
Rsn81_5 sn81_5 sn82_5 11.551961
Rsp81_6 sp81_6 sp82_6 11.551961
Rsn81_6 sn81_6 sn82_6 11.551961
Rsp81_7 sp81_7 sp82_7 11.551961
Rsn81_7 sn81_7 sn82_7 11.551961
Rsp81_8 sp81_8 sp82_8 11.551961
Rsn81_8 sn81_8 sn82_8 11.551961
Rsp81_9 sp81_9 sp82_9 11.551961
Rsn81_9 sn81_9 sn82_9 11.551961
Rsp81_10 sp81_10 sp82_10 11.551961
Rsn81_10 sn81_10 sn82_10 11.551961
Rsp81_11 sp81_11 sp82_11 11.551961
Rsn81_11 sn81_11 sn82_11 11.551961
Rsp81_12 sp81_12 sp82_12 11.551961
Rsn81_12 sn81_12 sn82_12 11.551961
Rsp81_13 sp81_13 sp82_13 11.551961
Rsn81_13 sn81_13 sn82_13 11.551961
Rsp81_14 sp81_14 sp82_14 11.551961
Rsn81_14 sn81_14 sn82_14 11.551961
Rsp81_15 sp81_15 sp82_15 11.551961
Rsn81_15 sn81_15 sn82_15 11.551961
Rsp81_16 sp81_16 sp82_16 11.551961
Rsn81_16 sn81_16 sn82_16 11.551961
Rsp81_17 sp81_17 sp82_17 11.551961
Rsn81_17 sn81_17 sn82_17 11.551961
Rsp81_18 sp81_18 sp82_18 11.551961
Rsn81_18 sn81_18 sn82_18 11.551961
Rsp81_19 sp81_19 sp82_19 11.551961
Rsn81_19 sn81_19 sn82_19 11.551961
Rsp81_20 sp81_20 sp82_20 11.551961
Rsn81_20 sn81_20 sn82_20 11.551961
Rsp81_21 sp81_21 sp82_21 11.551961
Rsn81_21 sn81_21 sn82_21 11.551961
Rsp81_22 sp81_22 sp82_22 11.551961
Rsn81_22 sn81_22 sn82_22 11.551961
Rsp81_23 sp81_23 sp82_23 11.551961
Rsn81_23 sn81_23 sn82_23 11.551961
Rsp81_24 sp81_24 sp82_24 11.551961
Rsn81_24 sn81_24 sn82_24 11.551961
Rsp81_25 sp81_25 sp82_25 11.551961
Rsn81_25 sn81_25 sn82_25 11.551961
Rsp81_26 sp81_26 sp82_26 11.551961
Rsn81_26 sn81_26 sn82_26 11.551961
Rsp81_27 sp81_27 sp82_27 11.551961
Rsn81_27 sn81_27 sn82_27 11.551961
Rsp81_28 sp81_28 sp82_28 11.551961
Rsn81_28 sn81_28 sn82_28 11.551961
Rsp81_29 sp81_29 sp82_29 11.551961
Rsn81_29 sn81_29 sn82_29 11.551961
Rsp81_30 sp81_30 sp82_30 11.551961
Rsn81_30 sn81_30 sn82_30 11.551961
Rsp81_31 sp81_31 sp82_31 11.551961
Rsn81_31 sn81_31 sn82_31 11.551961
Rsp81_32 sp81_32 sp82_32 11.551961
Rsn81_32 sn81_32 sn82_32 11.551961
Rsp81_33 sp81_33 sp82_33 11.551961
Rsn81_33 sn81_33 sn82_33 11.551961
Rsp81_34 sp81_34 sp82_34 11.551961
Rsn81_34 sn81_34 sn82_34 11.551961
Rsp81_35 sp81_35 sp82_35 11.551961
Rsn81_35 sn81_35 sn82_35 11.551961
Rsp81_36 sp81_36 sp82_36 11.551961
Rsn81_36 sn81_36 sn82_36 11.551961
Rsp81_37 sp81_37 sp82_37 11.551961
Rsn81_37 sn81_37 sn82_37 11.551961
Rsp81_38 sp81_38 sp82_38 11.551961
Rsn81_38 sn81_38 sn82_38 11.551961
Rsp81_39 sp81_39 sp82_39 11.551961
Rsn81_39 sn81_39 sn82_39 11.551961
Rsp81_40 sp81_40 sp82_40 11.551961
Rsn81_40 sn81_40 sn82_40 11.551961
Rsp81_41 sp81_41 sp82_41 11.551961
Rsn81_41 sn81_41 sn82_41 11.551961
Rsp81_42 sp81_42 sp82_42 11.551961
Rsn81_42 sn81_42 sn82_42 11.551961
Rsp81_43 sp81_43 sp82_43 11.551961
Rsn81_43 sn81_43 sn82_43 11.551961
Rsp81_44 sp81_44 sp82_44 11.551961
Rsn81_44 sn81_44 sn82_44 11.551961
Rsp81_45 sp81_45 sp82_45 11.551961
Rsn81_45 sn81_45 sn82_45 11.551961
Rsp81_46 sp81_46 sp82_46 11.551961
Rsn81_46 sn81_46 sn82_46 11.551961
Rsp81_47 sp81_47 sp82_47 11.551961
Rsn81_47 sn81_47 sn82_47 11.551961
Rsp81_48 sp81_48 sp82_48 11.551961
Rsn81_48 sn81_48 sn82_48 11.551961
Rsp81_49 sp81_49 sp82_49 11.551961
Rsn81_49 sn81_49 sn82_49 11.551961
Rsp81_50 sp81_50 sp82_50 11.551961
Rsn81_50 sn81_50 sn82_50 11.551961
Rsp81_51 sp81_51 sp82_51 11.551961
Rsn81_51 sn81_51 sn82_51 11.551961
Rsp81_52 sp81_52 sp82_52 11.551961
Rsn81_52 sn81_52 sn82_52 11.551961
Rsp81_53 sp81_53 sp82_53 11.551961
Rsn81_53 sn81_53 sn82_53 11.551961
Rsp81_54 sp81_54 sp82_54 11.551961
Rsn81_54 sn81_54 sn82_54 11.551961
Rsp81_55 sp81_55 sp82_55 11.551961
Rsn81_55 sn81_55 sn82_55 11.551961
Rsp81_56 sp81_56 sp82_56 11.551961
Rsn81_56 sn81_56 sn82_56 11.551961
Rsp81_57 sp81_57 sp82_57 11.551961
Rsn81_57 sn81_57 sn82_57 11.551961
Rsp81_58 sp81_58 sp82_58 11.551961
Rsn81_58 sn81_58 sn82_58 11.551961
Rsp81_59 sp81_59 sp82_59 11.551961
Rsn81_59 sn81_59 sn82_59 11.551961
Rsp81_60 sp81_60 sp82_60 11.551961
Rsn81_60 sn81_60 sn82_60 11.551961
Rsp81_61 sp81_61 sp82_61 11.551961
Rsn81_61 sn81_61 sn82_61 11.551961
Rsp81_62 sp81_62 sp82_62 11.551961
Rsn81_62 sn81_62 sn82_62 11.551961
Rsp81_63 sp81_63 sp82_63 11.551961
Rsn81_63 sn81_63 sn82_63 11.551961
Rsp81_64 sp81_64 sp82_64 11.551961
Rsn81_64 sn81_64 sn82_64 11.551961
Rsp81_65 sp81_65 sp82_65 11.551961
Rsn81_65 sn81_65 sn82_65 11.551961
Rsp81_66 sp81_66 sp82_66 11.551961
Rsn81_66 sn81_66 sn82_66 11.551961
Rsp81_67 sp81_67 sp82_67 11.551961
Rsn81_67 sn81_67 sn82_67 11.551961
Rsp81_68 sp81_68 sp82_68 11.551961
Rsn81_68 sn81_68 sn82_68 11.551961
Rsp81_69 sp81_69 sp82_69 11.551961
Rsn81_69 sn81_69 sn82_69 11.551961
Rsp81_70 sp81_70 sp82_70 11.551961
Rsn81_70 sn81_70 sn82_70 11.551961
Rsp81_71 sp81_71 sp82_71 11.551961
Rsn81_71 sn81_71 sn82_71 11.551961
Rsp81_72 sp81_72 sp82_72 11.551961
Rsn81_72 sn81_72 sn82_72 11.551961
Rsp81_73 sp81_73 sp82_73 11.551961
Rsn81_73 sn81_73 sn82_73 11.551961
Rsp81_74 sp81_74 sp82_74 11.551961
Rsn81_74 sn81_74 sn82_74 11.551961
Rsp81_75 sp81_75 sp82_75 11.551961
Rsn81_75 sn81_75 sn82_75 11.551961
Rsp81_76 sp81_76 sp82_76 11.551961
Rsn81_76 sn81_76 sn82_76 11.551961
Rsp81_77 sp81_77 sp82_77 11.551961
Rsn81_77 sn81_77 sn82_77 11.551961
Rsp81_78 sp81_78 sp82_78 11.551961
Rsn81_78 sn81_78 sn82_78 11.551961
Rsp81_79 sp81_79 sp82_79 11.551961
Rsn81_79 sn81_79 sn82_79 11.551961
Rsp81_80 sp81_80 sp82_80 11.551961
Rsn81_80 sn81_80 sn82_80 11.551961
Rsp81_81 sp81_81 sp82_81 11.551961
Rsn81_81 sn81_81 sn82_81 11.551961
Rsp81_82 sp81_82 sp82_82 11.551961
Rsn81_82 sn81_82 sn82_82 11.551961
Rsp81_83 sp81_83 sp82_83 11.551961
Rsn81_83 sn81_83 sn82_83 11.551961
Rsp81_84 sp81_84 sp82_84 11.551961
Rsn81_84 sn81_84 sn82_84 11.551961
Rsp82_1 sp82_1 sp83_1 11.551961
Rsn82_1 sn82_1 sn83_1 11.551961
Rsp82_2 sp82_2 sp83_2 11.551961
Rsn82_2 sn82_2 sn83_2 11.551961
Rsp82_3 sp82_3 sp83_3 11.551961
Rsn82_3 sn82_3 sn83_3 11.551961
Rsp82_4 sp82_4 sp83_4 11.551961
Rsn82_4 sn82_4 sn83_4 11.551961
Rsp82_5 sp82_5 sp83_5 11.551961
Rsn82_5 sn82_5 sn83_5 11.551961
Rsp82_6 sp82_6 sp83_6 11.551961
Rsn82_6 sn82_6 sn83_6 11.551961
Rsp82_7 sp82_7 sp83_7 11.551961
Rsn82_7 sn82_7 sn83_7 11.551961
Rsp82_8 sp82_8 sp83_8 11.551961
Rsn82_8 sn82_8 sn83_8 11.551961
Rsp82_9 sp82_9 sp83_9 11.551961
Rsn82_9 sn82_9 sn83_9 11.551961
Rsp82_10 sp82_10 sp83_10 11.551961
Rsn82_10 sn82_10 sn83_10 11.551961
Rsp82_11 sp82_11 sp83_11 11.551961
Rsn82_11 sn82_11 sn83_11 11.551961
Rsp82_12 sp82_12 sp83_12 11.551961
Rsn82_12 sn82_12 sn83_12 11.551961
Rsp82_13 sp82_13 sp83_13 11.551961
Rsn82_13 sn82_13 sn83_13 11.551961
Rsp82_14 sp82_14 sp83_14 11.551961
Rsn82_14 sn82_14 sn83_14 11.551961
Rsp82_15 sp82_15 sp83_15 11.551961
Rsn82_15 sn82_15 sn83_15 11.551961
Rsp82_16 sp82_16 sp83_16 11.551961
Rsn82_16 sn82_16 sn83_16 11.551961
Rsp82_17 sp82_17 sp83_17 11.551961
Rsn82_17 sn82_17 sn83_17 11.551961
Rsp82_18 sp82_18 sp83_18 11.551961
Rsn82_18 sn82_18 sn83_18 11.551961
Rsp82_19 sp82_19 sp83_19 11.551961
Rsn82_19 sn82_19 sn83_19 11.551961
Rsp82_20 sp82_20 sp83_20 11.551961
Rsn82_20 sn82_20 sn83_20 11.551961
Rsp82_21 sp82_21 sp83_21 11.551961
Rsn82_21 sn82_21 sn83_21 11.551961
Rsp82_22 sp82_22 sp83_22 11.551961
Rsn82_22 sn82_22 sn83_22 11.551961
Rsp82_23 sp82_23 sp83_23 11.551961
Rsn82_23 sn82_23 sn83_23 11.551961
Rsp82_24 sp82_24 sp83_24 11.551961
Rsn82_24 sn82_24 sn83_24 11.551961
Rsp82_25 sp82_25 sp83_25 11.551961
Rsn82_25 sn82_25 sn83_25 11.551961
Rsp82_26 sp82_26 sp83_26 11.551961
Rsn82_26 sn82_26 sn83_26 11.551961
Rsp82_27 sp82_27 sp83_27 11.551961
Rsn82_27 sn82_27 sn83_27 11.551961
Rsp82_28 sp82_28 sp83_28 11.551961
Rsn82_28 sn82_28 sn83_28 11.551961
Rsp82_29 sp82_29 sp83_29 11.551961
Rsn82_29 sn82_29 sn83_29 11.551961
Rsp82_30 sp82_30 sp83_30 11.551961
Rsn82_30 sn82_30 sn83_30 11.551961
Rsp82_31 sp82_31 sp83_31 11.551961
Rsn82_31 sn82_31 sn83_31 11.551961
Rsp82_32 sp82_32 sp83_32 11.551961
Rsn82_32 sn82_32 sn83_32 11.551961
Rsp82_33 sp82_33 sp83_33 11.551961
Rsn82_33 sn82_33 sn83_33 11.551961
Rsp82_34 sp82_34 sp83_34 11.551961
Rsn82_34 sn82_34 sn83_34 11.551961
Rsp82_35 sp82_35 sp83_35 11.551961
Rsn82_35 sn82_35 sn83_35 11.551961
Rsp82_36 sp82_36 sp83_36 11.551961
Rsn82_36 sn82_36 sn83_36 11.551961
Rsp82_37 sp82_37 sp83_37 11.551961
Rsn82_37 sn82_37 sn83_37 11.551961
Rsp82_38 sp82_38 sp83_38 11.551961
Rsn82_38 sn82_38 sn83_38 11.551961
Rsp82_39 sp82_39 sp83_39 11.551961
Rsn82_39 sn82_39 sn83_39 11.551961
Rsp82_40 sp82_40 sp83_40 11.551961
Rsn82_40 sn82_40 sn83_40 11.551961
Rsp82_41 sp82_41 sp83_41 11.551961
Rsn82_41 sn82_41 sn83_41 11.551961
Rsp82_42 sp82_42 sp83_42 11.551961
Rsn82_42 sn82_42 sn83_42 11.551961
Rsp82_43 sp82_43 sp83_43 11.551961
Rsn82_43 sn82_43 sn83_43 11.551961
Rsp82_44 sp82_44 sp83_44 11.551961
Rsn82_44 sn82_44 sn83_44 11.551961
Rsp82_45 sp82_45 sp83_45 11.551961
Rsn82_45 sn82_45 sn83_45 11.551961
Rsp82_46 sp82_46 sp83_46 11.551961
Rsn82_46 sn82_46 sn83_46 11.551961
Rsp82_47 sp82_47 sp83_47 11.551961
Rsn82_47 sn82_47 sn83_47 11.551961
Rsp82_48 sp82_48 sp83_48 11.551961
Rsn82_48 sn82_48 sn83_48 11.551961
Rsp82_49 sp82_49 sp83_49 11.551961
Rsn82_49 sn82_49 sn83_49 11.551961
Rsp82_50 sp82_50 sp83_50 11.551961
Rsn82_50 sn82_50 sn83_50 11.551961
Rsp82_51 sp82_51 sp83_51 11.551961
Rsn82_51 sn82_51 sn83_51 11.551961
Rsp82_52 sp82_52 sp83_52 11.551961
Rsn82_52 sn82_52 sn83_52 11.551961
Rsp82_53 sp82_53 sp83_53 11.551961
Rsn82_53 sn82_53 sn83_53 11.551961
Rsp82_54 sp82_54 sp83_54 11.551961
Rsn82_54 sn82_54 sn83_54 11.551961
Rsp82_55 sp82_55 sp83_55 11.551961
Rsn82_55 sn82_55 sn83_55 11.551961
Rsp82_56 sp82_56 sp83_56 11.551961
Rsn82_56 sn82_56 sn83_56 11.551961
Rsp82_57 sp82_57 sp83_57 11.551961
Rsn82_57 sn82_57 sn83_57 11.551961
Rsp82_58 sp82_58 sp83_58 11.551961
Rsn82_58 sn82_58 sn83_58 11.551961
Rsp82_59 sp82_59 sp83_59 11.551961
Rsn82_59 sn82_59 sn83_59 11.551961
Rsp82_60 sp82_60 sp83_60 11.551961
Rsn82_60 sn82_60 sn83_60 11.551961
Rsp82_61 sp82_61 sp83_61 11.551961
Rsn82_61 sn82_61 sn83_61 11.551961
Rsp82_62 sp82_62 sp83_62 11.551961
Rsn82_62 sn82_62 sn83_62 11.551961
Rsp82_63 sp82_63 sp83_63 11.551961
Rsn82_63 sn82_63 sn83_63 11.551961
Rsp82_64 sp82_64 sp83_64 11.551961
Rsn82_64 sn82_64 sn83_64 11.551961
Rsp82_65 sp82_65 sp83_65 11.551961
Rsn82_65 sn82_65 sn83_65 11.551961
Rsp82_66 sp82_66 sp83_66 11.551961
Rsn82_66 sn82_66 sn83_66 11.551961
Rsp82_67 sp82_67 sp83_67 11.551961
Rsn82_67 sn82_67 sn83_67 11.551961
Rsp82_68 sp82_68 sp83_68 11.551961
Rsn82_68 sn82_68 sn83_68 11.551961
Rsp82_69 sp82_69 sp83_69 11.551961
Rsn82_69 sn82_69 sn83_69 11.551961
Rsp82_70 sp82_70 sp83_70 11.551961
Rsn82_70 sn82_70 sn83_70 11.551961
Rsp82_71 sp82_71 sp83_71 11.551961
Rsn82_71 sn82_71 sn83_71 11.551961
Rsp82_72 sp82_72 sp83_72 11.551961
Rsn82_72 sn82_72 sn83_72 11.551961
Rsp82_73 sp82_73 sp83_73 11.551961
Rsn82_73 sn82_73 sn83_73 11.551961
Rsp82_74 sp82_74 sp83_74 11.551961
Rsn82_74 sn82_74 sn83_74 11.551961
Rsp82_75 sp82_75 sp83_75 11.551961
Rsn82_75 sn82_75 sn83_75 11.551961
Rsp82_76 sp82_76 sp83_76 11.551961
Rsn82_76 sn82_76 sn83_76 11.551961
Rsp82_77 sp82_77 sp83_77 11.551961
Rsn82_77 sn82_77 sn83_77 11.551961
Rsp82_78 sp82_78 sp83_78 11.551961
Rsn82_78 sn82_78 sn83_78 11.551961
Rsp82_79 sp82_79 sp83_79 11.551961
Rsn82_79 sn82_79 sn83_79 11.551961
Rsp82_80 sp82_80 sp83_80 11.551961
Rsn82_80 sn82_80 sn83_80 11.551961
Rsp82_81 sp82_81 sp83_81 11.551961
Rsn82_81 sn82_81 sn83_81 11.551961
Rsp82_82 sp82_82 sp83_82 11.551961
Rsn82_82 sn82_82 sn83_82 11.551961
Rsp82_83 sp82_83 sp83_83 11.551961
Rsn82_83 sn82_83 sn83_83 11.551961
Rsp82_84 sp82_84 sp83_84 11.551961
Rsn82_84 sn82_84 sn83_84 11.551961
Rsp83_1 sp83_1 sp84_1 11.551961
Rsn83_1 sn83_1 sn84_1 11.551961
Rsp83_2 sp83_2 sp84_2 11.551961
Rsn83_2 sn83_2 sn84_2 11.551961
Rsp83_3 sp83_3 sp84_3 11.551961
Rsn83_3 sn83_3 sn84_3 11.551961
Rsp83_4 sp83_4 sp84_4 11.551961
Rsn83_4 sn83_4 sn84_4 11.551961
Rsp83_5 sp83_5 sp84_5 11.551961
Rsn83_5 sn83_5 sn84_5 11.551961
Rsp83_6 sp83_6 sp84_6 11.551961
Rsn83_6 sn83_6 sn84_6 11.551961
Rsp83_7 sp83_7 sp84_7 11.551961
Rsn83_7 sn83_7 sn84_7 11.551961
Rsp83_8 sp83_8 sp84_8 11.551961
Rsn83_8 sn83_8 sn84_8 11.551961
Rsp83_9 sp83_9 sp84_9 11.551961
Rsn83_9 sn83_9 sn84_9 11.551961
Rsp83_10 sp83_10 sp84_10 11.551961
Rsn83_10 sn83_10 sn84_10 11.551961
Rsp83_11 sp83_11 sp84_11 11.551961
Rsn83_11 sn83_11 sn84_11 11.551961
Rsp83_12 sp83_12 sp84_12 11.551961
Rsn83_12 sn83_12 sn84_12 11.551961
Rsp83_13 sp83_13 sp84_13 11.551961
Rsn83_13 sn83_13 sn84_13 11.551961
Rsp83_14 sp83_14 sp84_14 11.551961
Rsn83_14 sn83_14 sn84_14 11.551961
Rsp83_15 sp83_15 sp84_15 11.551961
Rsn83_15 sn83_15 sn84_15 11.551961
Rsp83_16 sp83_16 sp84_16 11.551961
Rsn83_16 sn83_16 sn84_16 11.551961
Rsp83_17 sp83_17 sp84_17 11.551961
Rsn83_17 sn83_17 sn84_17 11.551961
Rsp83_18 sp83_18 sp84_18 11.551961
Rsn83_18 sn83_18 sn84_18 11.551961
Rsp83_19 sp83_19 sp84_19 11.551961
Rsn83_19 sn83_19 sn84_19 11.551961
Rsp83_20 sp83_20 sp84_20 11.551961
Rsn83_20 sn83_20 sn84_20 11.551961
Rsp83_21 sp83_21 sp84_21 11.551961
Rsn83_21 sn83_21 sn84_21 11.551961
Rsp83_22 sp83_22 sp84_22 11.551961
Rsn83_22 sn83_22 sn84_22 11.551961
Rsp83_23 sp83_23 sp84_23 11.551961
Rsn83_23 sn83_23 sn84_23 11.551961
Rsp83_24 sp83_24 sp84_24 11.551961
Rsn83_24 sn83_24 sn84_24 11.551961
Rsp83_25 sp83_25 sp84_25 11.551961
Rsn83_25 sn83_25 sn84_25 11.551961
Rsp83_26 sp83_26 sp84_26 11.551961
Rsn83_26 sn83_26 sn84_26 11.551961
Rsp83_27 sp83_27 sp84_27 11.551961
Rsn83_27 sn83_27 sn84_27 11.551961
Rsp83_28 sp83_28 sp84_28 11.551961
Rsn83_28 sn83_28 sn84_28 11.551961
Rsp83_29 sp83_29 sp84_29 11.551961
Rsn83_29 sn83_29 sn84_29 11.551961
Rsp83_30 sp83_30 sp84_30 11.551961
Rsn83_30 sn83_30 sn84_30 11.551961
Rsp83_31 sp83_31 sp84_31 11.551961
Rsn83_31 sn83_31 sn84_31 11.551961
Rsp83_32 sp83_32 sp84_32 11.551961
Rsn83_32 sn83_32 sn84_32 11.551961
Rsp83_33 sp83_33 sp84_33 11.551961
Rsn83_33 sn83_33 sn84_33 11.551961
Rsp83_34 sp83_34 sp84_34 11.551961
Rsn83_34 sn83_34 sn84_34 11.551961
Rsp83_35 sp83_35 sp84_35 11.551961
Rsn83_35 sn83_35 sn84_35 11.551961
Rsp83_36 sp83_36 sp84_36 11.551961
Rsn83_36 sn83_36 sn84_36 11.551961
Rsp83_37 sp83_37 sp84_37 11.551961
Rsn83_37 sn83_37 sn84_37 11.551961
Rsp83_38 sp83_38 sp84_38 11.551961
Rsn83_38 sn83_38 sn84_38 11.551961
Rsp83_39 sp83_39 sp84_39 11.551961
Rsn83_39 sn83_39 sn84_39 11.551961
Rsp83_40 sp83_40 sp84_40 11.551961
Rsn83_40 sn83_40 sn84_40 11.551961
Rsp83_41 sp83_41 sp84_41 11.551961
Rsn83_41 sn83_41 sn84_41 11.551961
Rsp83_42 sp83_42 sp84_42 11.551961
Rsn83_42 sn83_42 sn84_42 11.551961
Rsp83_43 sp83_43 sp84_43 11.551961
Rsn83_43 sn83_43 sn84_43 11.551961
Rsp83_44 sp83_44 sp84_44 11.551961
Rsn83_44 sn83_44 sn84_44 11.551961
Rsp83_45 sp83_45 sp84_45 11.551961
Rsn83_45 sn83_45 sn84_45 11.551961
Rsp83_46 sp83_46 sp84_46 11.551961
Rsn83_46 sn83_46 sn84_46 11.551961
Rsp83_47 sp83_47 sp84_47 11.551961
Rsn83_47 sn83_47 sn84_47 11.551961
Rsp83_48 sp83_48 sp84_48 11.551961
Rsn83_48 sn83_48 sn84_48 11.551961
Rsp83_49 sp83_49 sp84_49 11.551961
Rsn83_49 sn83_49 sn84_49 11.551961
Rsp83_50 sp83_50 sp84_50 11.551961
Rsn83_50 sn83_50 sn84_50 11.551961
Rsp83_51 sp83_51 sp84_51 11.551961
Rsn83_51 sn83_51 sn84_51 11.551961
Rsp83_52 sp83_52 sp84_52 11.551961
Rsn83_52 sn83_52 sn84_52 11.551961
Rsp83_53 sp83_53 sp84_53 11.551961
Rsn83_53 sn83_53 sn84_53 11.551961
Rsp83_54 sp83_54 sp84_54 11.551961
Rsn83_54 sn83_54 sn84_54 11.551961
Rsp83_55 sp83_55 sp84_55 11.551961
Rsn83_55 sn83_55 sn84_55 11.551961
Rsp83_56 sp83_56 sp84_56 11.551961
Rsn83_56 sn83_56 sn84_56 11.551961
Rsp83_57 sp83_57 sp84_57 11.551961
Rsn83_57 sn83_57 sn84_57 11.551961
Rsp83_58 sp83_58 sp84_58 11.551961
Rsn83_58 sn83_58 sn84_58 11.551961
Rsp83_59 sp83_59 sp84_59 11.551961
Rsn83_59 sn83_59 sn84_59 11.551961
Rsp83_60 sp83_60 sp84_60 11.551961
Rsn83_60 sn83_60 sn84_60 11.551961
Rsp83_61 sp83_61 sp84_61 11.551961
Rsn83_61 sn83_61 sn84_61 11.551961
Rsp83_62 sp83_62 sp84_62 11.551961
Rsn83_62 sn83_62 sn84_62 11.551961
Rsp83_63 sp83_63 sp84_63 11.551961
Rsn83_63 sn83_63 sn84_63 11.551961
Rsp83_64 sp83_64 sp84_64 11.551961
Rsn83_64 sn83_64 sn84_64 11.551961
Rsp83_65 sp83_65 sp84_65 11.551961
Rsn83_65 sn83_65 sn84_65 11.551961
Rsp83_66 sp83_66 sp84_66 11.551961
Rsn83_66 sn83_66 sn84_66 11.551961
Rsp83_67 sp83_67 sp84_67 11.551961
Rsn83_67 sn83_67 sn84_67 11.551961
Rsp83_68 sp83_68 sp84_68 11.551961
Rsn83_68 sn83_68 sn84_68 11.551961
Rsp83_69 sp83_69 sp84_69 11.551961
Rsn83_69 sn83_69 sn84_69 11.551961
Rsp83_70 sp83_70 sp84_70 11.551961
Rsn83_70 sn83_70 sn84_70 11.551961
Rsp83_71 sp83_71 sp84_71 11.551961
Rsn83_71 sn83_71 sn84_71 11.551961
Rsp83_72 sp83_72 sp84_72 11.551961
Rsn83_72 sn83_72 sn84_72 11.551961
Rsp83_73 sp83_73 sp84_73 11.551961
Rsn83_73 sn83_73 sn84_73 11.551961
Rsp83_74 sp83_74 sp84_74 11.551961
Rsn83_74 sn83_74 sn84_74 11.551961
Rsp83_75 sp83_75 sp84_75 11.551961
Rsn83_75 sn83_75 sn84_75 11.551961
Rsp83_76 sp83_76 sp84_76 11.551961
Rsn83_76 sn83_76 sn84_76 11.551961
Rsp83_77 sp83_77 sp84_77 11.551961
Rsn83_77 sn83_77 sn84_77 11.551961
Rsp83_78 sp83_78 sp84_78 11.551961
Rsn83_78 sn83_78 sn84_78 11.551961
Rsp83_79 sp83_79 sp84_79 11.551961
Rsn83_79 sn83_79 sn84_79 11.551961
Rsp83_80 sp83_80 sp84_80 11.551961
Rsn83_80 sn83_80 sn84_80 11.551961
Rsp83_81 sp83_81 sp84_81 11.551961
Rsn83_81 sn83_81 sn84_81 11.551961
Rsp83_82 sp83_82 sp84_82 11.551961
Rsn83_82 sn83_82 sn84_82 11.551961
Rsp83_83 sp83_83 sp84_83 11.551961
Rsn83_83 sn83_83 sn84_83 11.551961
Rsp83_84 sp83_84 sp84_84 11.551961
Rsn83_84 sn83_84 sn84_84 11.551961
Rsp84_1 sp84_1 sp85_1 11.551961
Rsn84_1 sn84_1 sn85_1 11.551961
Rsp84_2 sp84_2 sp85_2 11.551961
Rsn84_2 sn84_2 sn85_2 11.551961
Rsp84_3 sp84_3 sp85_3 11.551961
Rsn84_3 sn84_3 sn85_3 11.551961
Rsp84_4 sp84_4 sp85_4 11.551961
Rsn84_4 sn84_4 sn85_4 11.551961
Rsp84_5 sp84_5 sp85_5 11.551961
Rsn84_5 sn84_5 sn85_5 11.551961
Rsp84_6 sp84_6 sp85_6 11.551961
Rsn84_6 sn84_6 sn85_6 11.551961
Rsp84_7 sp84_7 sp85_7 11.551961
Rsn84_7 sn84_7 sn85_7 11.551961
Rsp84_8 sp84_8 sp85_8 11.551961
Rsn84_8 sn84_8 sn85_8 11.551961
Rsp84_9 sp84_9 sp85_9 11.551961
Rsn84_9 sn84_9 sn85_9 11.551961
Rsp84_10 sp84_10 sp85_10 11.551961
Rsn84_10 sn84_10 sn85_10 11.551961
Rsp84_11 sp84_11 sp85_11 11.551961
Rsn84_11 sn84_11 sn85_11 11.551961
Rsp84_12 sp84_12 sp85_12 11.551961
Rsn84_12 sn84_12 sn85_12 11.551961
Rsp84_13 sp84_13 sp85_13 11.551961
Rsn84_13 sn84_13 sn85_13 11.551961
Rsp84_14 sp84_14 sp85_14 11.551961
Rsn84_14 sn84_14 sn85_14 11.551961
Rsp84_15 sp84_15 sp85_15 11.551961
Rsn84_15 sn84_15 sn85_15 11.551961
Rsp84_16 sp84_16 sp85_16 11.551961
Rsn84_16 sn84_16 sn85_16 11.551961
Rsp84_17 sp84_17 sp85_17 11.551961
Rsn84_17 sn84_17 sn85_17 11.551961
Rsp84_18 sp84_18 sp85_18 11.551961
Rsn84_18 sn84_18 sn85_18 11.551961
Rsp84_19 sp84_19 sp85_19 11.551961
Rsn84_19 sn84_19 sn85_19 11.551961
Rsp84_20 sp84_20 sp85_20 11.551961
Rsn84_20 sn84_20 sn85_20 11.551961
Rsp84_21 sp84_21 sp85_21 11.551961
Rsn84_21 sn84_21 sn85_21 11.551961
Rsp84_22 sp84_22 sp85_22 11.551961
Rsn84_22 sn84_22 sn85_22 11.551961
Rsp84_23 sp84_23 sp85_23 11.551961
Rsn84_23 sn84_23 sn85_23 11.551961
Rsp84_24 sp84_24 sp85_24 11.551961
Rsn84_24 sn84_24 sn85_24 11.551961
Rsp84_25 sp84_25 sp85_25 11.551961
Rsn84_25 sn84_25 sn85_25 11.551961
Rsp84_26 sp84_26 sp85_26 11.551961
Rsn84_26 sn84_26 sn85_26 11.551961
Rsp84_27 sp84_27 sp85_27 11.551961
Rsn84_27 sn84_27 sn85_27 11.551961
Rsp84_28 sp84_28 sp85_28 11.551961
Rsn84_28 sn84_28 sn85_28 11.551961
Rsp84_29 sp84_29 sp85_29 11.551961
Rsn84_29 sn84_29 sn85_29 11.551961
Rsp84_30 sp84_30 sp85_30 11.551961
Rsn84_30 sn84_30 sn85_30 11.551961
Rsp84_31 sp84_31 sp85_31 11.551961
Rsn84_31 sn84_31 sn85_31 11.551961
Rsp84_32 sp84_32 sp85_32 11.551961
Rsn84_32 sn84_32 sn85_32 11.551961
Rsp84_33 sp84_33 sp85_33 11.551961
Rsn84_33 sn84_33 sn85_33 11.551961
Rsp84_34 sp84_34 sp85_34 11.551961
Rsn84_34 sn84_34 sn85_34 11.551961
Rsp84_35 sp84_35 sp85_35 11.551961
Rsn84_35 sn84_35 sn85_35 11.551961
Rsp84_36 sp84_36 sp85_36 11.551961
Rsn84_36 sn84_36 sn85_36 11.551961
Rsp84_37 sp84_37 sp85_37 11.551961
Rsn84_37 sn84_37 sn85_37 11.551961
Rsp84_38 sp84_38 sp85_38 11.551961
Rsn84_38 sn84_38 sn85_38 11.551961
Rsp84_39 sp84_39 sp85_39 11.551961
Rsn84_39 sn84_39 sn85_39 11.551961
Rsp84_40 sp84_40 sp85_40 11.551961
Rsn84_40 sn84_40 sn85_40 11.551961
Rsp84_41 sp84_41 sp85_41 11.551961
Rsn84_41 sn84_41 sn85_41 11.551961
Rsp84_42 sp84_42 sp85_42 11.551961
Rsn84_42 sn84_42 sn85_42 11.551961
Rsp84_43 sp84_43 sp85_43 11.551961
Rsn84_43 sn84_43 sn85_43 11.551961
Rsp84_44 sp84_44 sp85_44 11.551961
Rsn84_44 sn84_44 sn85_44 11.551961
Rsp84_45 sp84_45 sp85_45 11.551961
Rsn84_45 sn84_45 sn85_45 11.551961
Rsp84_46 sp84_46 sp85_46 11.551961
Rsn84_46 sn84_46 sn85_46 11.551961
Rsp84_47 sp84_47 sp85_47 11.551961
Rsn84_47 sn84_47 sn85_47 11.551961
Rsp84_48 sp84_48 sp85_48 11.551961
Rsn84_48 sn84_48 sn85_48 11.551961
Rsp84_49 sp84_49 sp85_49 11.551961
Rsn84_49 sn84_49 sn85_49 11.551961
Rsp84_50 sp84_50 sp85_50 11.551961
Rsn84_50 sn84_50 sn85_50 11.551961
Rsp84_51 sp84_51 sp85_51 11.551961
Rsn84_51 sn84_51 sn85_51 11.551961
Rsp84_52 sp84_52 sp85_52 11.551961
Rsn84_52 sn84_52 sn85_52 11.551961
Rsp84_53 sp84_53 sp85_53 11.551961
Rsn84_53 sn84_53 sn85_53 11.551961
Rsp84_54 sp84_54 sp85_54 11.551961
Rsn84_54 sn84_54 sn85_54 11.551961
Rsp84_55 sp84_55 sp85_55 11.551961
Rsn84_55 sn84_55 sn85_55 11.551961
Rsp84_56 sp84_56 sp85_56 11.551961
Rsn84_56 sn84_56 sn85_56 11.551961
Rsp84_57 sp84_57 sp85_57 11.551961
Rsn84_57 sn84_57 sn85_57 11.551961
Rsp84_58 sp84_58 sp85_58 11.551961
Rsn84_58 sn84_58 sn85_58 11.551961
Rsp84_59 sp84_59 sp85_59 11.551961
Rsn84_59 sn84_59 sn85_59 11.551961
Rsp84_60 sp84_60 sp85_60 11.551961
Rsn84_60 sn84_60 sn85_60 11.551961
Rsp84_61 sp84_61 sp85_61 11.551961
Rsn84_61 sn84_61 sn85_61 11.551961
Rsp84_62 sp84_62 sp85_62 11.551961
Rsn84_62 sn84_62 sn85_62 11.551961
Rsp84_63 sp84_63 sp85_63 11.551961
Rsn84_63 sn84_63 sn85_63 11.551961
Rsp84_64 sp84_64 sp85_64 11.551961
Rsn84_64 sn84_64 sn85_64 11.551961
Rsp84_65 sp84_65 sp85_65 11.551961
Rsn84_65 sn84_65 sn85_65 11.551961
Rsp84_66 sp84_66 sp85_66 11.551961
Rsn84_66 sn84_66 sn85_66 11.551961
Rsp84_67 sp84_67 sp85_67 11.551961
Rsn84_67 sn84_67 sn85_67 11.551961
Rsp84_68 sp84_68 sp85_68 11.551961
Rsn84_68 sn84_68 sn85_68 11.551961
Rsp84_69 sp84_69 sp85_69 11.551961
Rsn84_69 sn84_69 sn85_69 11.551961
Rsp84_70 sp84_70 sp85_70 11.551961
Rsn84_70 sn84_70 sn85_70 11.551961
Rsp84_71 sp84_71 sp85_71 11.551961
Rsn84_71 sn84_71 sn85_71 11.551961
Rsp84_72 sp84_72 sp85_72 11.551961
Rsn84_72 sn84_72 sn85_72 11.551961
Rsp84_73 sp84_73 sp85_73 11.551961
Rsn84_73 sn84_73 sn85_73 11.551961
Rsp84_74 sp84_74 sp85_74 11.551961
Rsn84_74 sn84_74 sn85_74 11.551961
Rsp84_75 sp84_75 sp85_75 11.551961
Rsn84_75 sn84_75 sn85_75 11.551961
Rsp84_76 sp84_76 sp85_76 11.551961
Rsn84_76 sn84_76 sn85_76 11.551961
Rsp84_77 sp84_77 sp85_77 11.551961
Rsn84_77 sn84_77 sn85_77 11.551961
Rsp84_78 sp84_78 sp85_78 11.551961
Rsn84_78 sn84_78 sn85_78 11.551961
Rsp84_79 sp84_79 sp85_79 11.551961
Rsn84_79 sn84_79 sn85_79 11.551961
Rsp84_80 sp84_80 sp85_80 11.551961
Rsn84_80 sn84_80 sn85_80 11.551961
Rsp84_81 sp84_81 sp85_81 11.551961
Rsn84_81 sn84_81 sn85_81 11.551961
Rsp84_82 sp84_82 sp85_82 11.551961
Rsn84_82 sn84_82 sn85_82 11.551961
Rsp84_83 sp84_83 sp85_83 11.551961
Rsn84_83 sn84_83 sn85_83 11.551961
Rsp84_84 sp84_84 sp85_84 11.551961
Rsn84_84 sn84_84 sn85_84 11.551961
Rsp85_1 sp85_1 sp86_1 11.551961
Rsn85_1 sn85_1 sn86_1 11.551961
Rsp85_2 sp85_2 sp86_2 11.551961
Rsn85_2 sn85_2 sn86_2 11.551961
Rsp85_3 sp85_3 sp86_3 11.551961
Rsn85_3 sn85_3 sn86_3 11.551961
Rsp85_4 sp85_4 sp86_4 11.551961
Rsn85_4 sn85_4 sn86_4 11.551961
Rsp85_5 sp85_5 sp86_5 11.551961
Rsn85_5 sn85_5 sn86_5 11.551961
Rsp85_6 sp85_6 sp86_6 11.551961
Rsn85_6 sn85_6 sn86_6 11.551961
Rsp85_7 sp85_7 sp86_7 11.551961
Rsn85_7 sn85_7 sn86_7 11.551961
Rsp85_8 sp85_8 sp86_8 11.551961
Rsn85_8 sn85_8 sn86_8 11.551961
Rsp85_9 sp85_9 sp86_9 11.551961
Rsn85_9 sn85_9 sn86_9 11.551961
Rsp85_10 sp85_10 sp86_10 11.551961
Rsn85_10 sn85_10 sn86_10 11.551961
Rsp85_11 sp85_11 sp86_11 11.551961
Rsn85_11 sn85_11 sn86_11 11.551961
Rsp85_12 sp85_12 sp86_12 11.551961
Rsn85_12 sn85_12 sn86_12 11.551961
Rsp85_13 sp85_13 sp86_13 11.551961
Rsn85_13 sn85_13 sn86_13 11.551961
Rsp85_14 sp85_14 sp86_14 11.551961
Rsn85_14 sn85_14 sn86_14 11.551961
Rsp85_15 sp85_15 sp86_15 11.551961
Rsn85_15 sn85_15 sn86_15 11.551961
Rsp85_16 sp85_16 sp86_16 11.551961
Rsn85_16 sn85_16 sn86_16 11.551961
Rsp85_17 sp85_17 sp86_17 11.551961
Rsn85_17 sn85_17 sn86_17 11.551961
Rsp85_18 sp85_18 sp86_18 11.551961
Rsn85_18 sn85_18 sn86_18 11.551961
Rsp85_19 sp85_19 sp86_19 11.551961
Rsn85_19 sn85_19 sn86_19 11.551961
Rsp85_20 sp85_20 sp86_20 11.551961
Rsn85_20 sn85_20 sn86_20 11.551961
Rsp85_21 sp85_21 sp86_21 11.551961
Rsn85_21 sn85_21 sn86_21 11.551961
Rsp85_22 sp85_22 sp86_22 11.551961
Rsn85_22 sn85_22 sn86_22 11.551961
Rsp85_23 sp85_23 sp86_23 11.551961
Rsn85_23 sn85_23 sn86_23 11.551961
Rsp85_24 sp85_24 sp86_24 11.551961
Rsn85_24 sn85_24 sn86_24 11.551961
Rsp85_25 sp85_25 sp86_25 11.551961
Rsn85_25 sn85_25 sn86_25 11.551961
Rsp85_26 sp85_26 sp86_26 11.551961
Rsn85_26 sn85_26 sn86_26 11.551961
Rsp85_27 sp85_27 sp86_27 11.551961
Rsn85_27 sn85_27 sn86_27 11.551961
Rsp85_28 sp85_28 sp86_28 11.551961
Rsn85_28 sn85_28 sn86_28 11.551961
Rsp85_29 sp85_29 sp86_29 11.551961
Rsn85_29 sn85_29 sn86_29 11.551961
Rsp85_30 sp85_30 sp86_30 11.551961
Rsn85_30 sn85_30 sn86_30 11.551961
Rsp85_31 sp85_31 sp86_31 11.551961
Rsn85_31 sn85_31 sn86_31 11.551961
Rsp85_32 sp85_32 sp86_32 11.551961
Rsn85_32 sn85_32 sn86_32 11.551961
Rsp85_33 sp85_33 sp86_33 11.551961
Rsn85_33 sn85_33 sn86_33 11.551961
Rsp85_34 sp85_34 sp86_34 11.551961
Rsn85_34 sn85_34 sn86_34 11.551961
Rsp85_35 sp85_35 sp86_35 11.551961
Rsn85_35 sn85_35 sn86_35 11.551961
Rsp85_36 sp85_36 sp86_36 11.551961
Rsn85_36 sn85_36 sn86_36 11.551961
Rsp85_37 sp85_37 sp86_37 11.551961
Rsn85_37 sn85_37 sn86_37 11.551961
Rsp85_38 sp85_38 sp86_38 11.551961
Rsn85_38 sn85_38 sn86_38 11.551961
Rsp85_39 sp85_39 sp86_39 11.551961
Rsn85_39 sn85_39 sn86_39 11.551961
Rsp85_40 sp85_40 sp86_40 11.551961
Rsn85_40 sn85_40 sn86_40 11.551961
Rsp85_41 sp85_41 sp86_41 11.551961
Rsn85_41 sn85_41 sn86_41 11.551961
Rsp85_42 sp85_42 sp86_42 11.551961
Rsn85_42 sn85_42 sn86_42 11.551961
Rsp85_43 sp85_43 sp86_43 11.551961
Rsn85_43 sn85_43 sn86_43 11.551961
Rsp85_44 sp85_44 sp86_44 11.551961
Rsn85_44 sn85_44 sn86_44 11.551961
Rsp85_45 sp85_45 sp86_45 11.551961
Rsn85_45 sn85_45 sn86_45 11.551961
Rsp85_46 sp85_46 sp86_46 11.551961
Rsn85_46 sn85_46 sn86_46 11.551961
Rsp85_47 sp85_47 sp86_47 11.551961
Rsn85_47 sn85_47 sn86_47 11.551961
Rsp85_48 sp85_48 sp86_48 11.551961
Rsn85_48 sn85_48 sn86_48 11.551961
Rsp85_49 sp85_49 sp86_49 11.551961
Rsn85_49 sn85_49 sn86_49 11.551961
Rsp85_50 sp85_50 sp86_50 11.551961
Rsn85_50 sn85_50 sn86_50 11.551961
Rsp85_51 sp85_51 sp86_51 11.551961
Rsn85_51 sn85_51 sn86_51 11.551961
Rsp85_52 sp85_52 sp86_52 11.551961
Rsn85_52 sn85_52 sn86_52 11.551961
Rsp85_53 sp85_53 sp86_53 11.551961
Rsn85_53 sn85_53 sn86_53 11.551961
Rsp85_54 sp85_54 sp86_54 11.551961
Rsn85_54 sn85_54 sn86_54 11.551961
Rsp85_55 sp85_55 sp86_55 11.551961
Rsn85_55 sn85_55 sn86_55 11.551961
Rsp85_56 sp85_56 sp86_56 11.551961
Rsn85_56 sn85_56 sn86_56 11.551961
Rsp85_57 sp85_57 sp86_57 11.551961
Rsn85_57 sn85_57 sn86_57 11.551961
Rsp85_58 sp85_58 sp86_58 11.551961
Rsn85_58 sn85_58 sn86_58 11.551961
Rsp85_59 sp85_59 sp86_59 11.551961
Rsn85_59 sn85_59 sn86_59 11.551961
Rsp85_60 sp85_60 sp86_60 11.551961
Rsn85_60 sn85_60 sn86_60 11.551961
Rsp85_61 sp85_61 sp86_61 11.551961
Rsn85_61 sn85_61 sn86_61 11.551961
Rsp85_62 sp85_62 sp86_62 11.551961
Rsn85_62 sn85_62 sn86_62 11.551961
Rsp85_63 sp85_63 sp86_63 11.551961
Rsn85_63 sn85_63 sn86_63 11.551961
Rsp85_64 sp85_64 sp86_64 11.551961
Rsn85_64 sn85_64 sn86_64 11.551961
Rsp85_65 sp85_65 sp86_65 11.551961
Rsn85_65 sn85_65 sn86_65 11.551961
Rsp85_66 sp85_66 sp86_66 11.551961
Rsn85_66 sn85_66 sn86_66 11.551961
Rsp85_67 sp85_67 sp86_67 11.551961
Rsn85_67 sn85_67 sn86_67 11.551961
Rsp85_68 sp85_68 sp86_68 11.551961
Rsn85_68 sn85_68 sn86_68 11.551961
Rsp85_69 sp85_69 sp86_69 11.551961
Rsn85_69 sn85_69 sn86_69 11.551961
Rsp85_70 sp85_70 sp86_70 11.551961
Rsn85_70 sn85_70 sn86_70 11.551961
Rsp85_71 sp85_71 sp86_71 11.551961
Rsn85_71 sn85_71 sn86_71 11.551961
Rsp85_72 sp85_72 sp86_72 11.551961
Rsn85_72 sn85_72 sn86_72 11.551961
Rsp85_73 sp85_73 sp86_73 11.551961
Rsn85_73 sn85_73 sn86_73 11.551961
Rsp85_74 sp85_74 sp86_74 11.551961
Rsn85_74 sn85_74 sn86_74 11.551961
Rsp85_75 sp85_75 sp86_75 11.551961
Rsn85_75 sn85_75 sn86_75 11.551961
Rsp85_76 sp85_76 sp86_76 11.551961
Rsn85_76 sn85_76 sn86_76 11.551961
Rsp85_77 sp85_77 sp86_77 11.551961
Rsn85_77 sn85_77 sn86_77 11.551961
Rsp85_78 sp85_78 sp86_78 11.551961
Rsn85_78 sn85_78 sn86_78 11.551961
Rsp85_79 sp85_79 sp86_79 11.551961
Rsn85_79 sn85_79 sn86_79 11.551961
Rsp85_80 sp85_80 sp86_80 11.551961
Rsn85_80 sn85_80 sn86_80 11.551961
Rsp85_81 sp85_81 sp86_81 11.551961
Rsn85_81 sn85_81 sn86_81 11.551961
Rsp85_82 sp85_82 sp86_82 11.551961
Rsn85_82 sn85_82 sn86_82 11.551961
Rsp85_83 sp85_83 sp86_83 11.551961
Rsn85_83 sn85_83 sn86_83 11.551961
Rsp85_84 sp85_84 sp86_84 11.551961
Rsn85_84 sn85_84 sn86_84 11.551961
Rsp86_1 sp86_1 sp87_1 11.551961
Rsn86_1 sn86_1 sn87_1 11.551961
Rsp86_2 sp86_2 sp87_2 11.551961
Rsn86_2 sn86_2 sn87_2 11.551961
Rsp86_3 sp86_3 sp87_3 11.551961
Rsn86_3 sn86_3 sn87_3 11.551961
Rsp86_4 sp86_4 sp87_4 11.551961
Rsn86_4 sn86_4 sn87_4 11.551961
Rsp86_5 sp86_5 sp87_5 11.551961
Rsn86_5 sn86_5 sn87_5 11.551961
Rsp86_6 sp86_6 sp87_6 11.551961
Rsn86_6 sn86_6 sn87_6 11.551961
Rsp86_7 sp86_7 sp87_7 11.551961
Rsn86_7 sn86_7 sn87_7 11.551961
Rsp86_8 sp86_8 sp87_8 11.551961
Rsn86_8 sn86_8 sn87_8 11.551961
Rsp86_9 sp86_9 sp87_9 11.551961
Rsn86_9 sn86_9 sn87_9 11.551961
Rsp86_10 sp86_10 sp87_10 11.551961
Rsn86_10 sn86_10 sn87_10 11.551961
Rsp86_11 sp86_11 sp87_11 11.551961
Rsn86_11 sn86_11 sn87_11 11.551961
Rsp86_12 sp86_12 sp87_12 11.551961
Rsn86_12 sn86_12 sn87_12 11.551961
Rsp86_13 sp86_13 sp87_13 11.551961
Rsn86_13 sn86_13 sn87_13 11.551961
Rsp86_14 sp86_14 sp87_14 11.551961
Rsn86_14 sn86_14 sn87_14 11.551961
Rsp86_15 sp86_15 sp87_15 11.551961
Rsn86_15 sn86_15 sn87_15 11.551961
Rsp86_16 sp86_16 sp87_16 11.551961
Rsn86_16 sn86_16 sn87_16 11.551961
Rsp86_17 sp86_17 sp87_17 11.551961
Rsn86_17 sn86_17 sn87_17 11.551961
Rsp86_18 sp86_18 sp87_18 11.551961
Rsn86_18 sn86_18 sn87_18 11.551961
Rsp86_19 sp86_19 sp87_19 11.551961
Rsn86_19 sn86_19 sn87_19 11.551961
Rsp86_20 sp86_20 sp87_20 11.551961
Rsn86_20 sn86_20 sn87_20 11.551961
Rsp86_21 sp86_21 sp87_21 11.551961
Rsn86_21 sn86_21 sn87_21 11.551961
Rsp86_22 sp86_22 sp87_22 11.551961
Rsn86_22 sn86_22 sn87_22 11.551961
Rsp86_23 sp86_23 sp87_23 11.551961
Rsn86_23 sn86_23 sn87_23 11.551961
Rsp86_24 sp86_24 sp87_24 11.551961
Rsn86_24 sn86_24 sn87_24 11.551961
Rsp86_25 sp86_25 sp87_25 11.551961
Rsn86_25 sn86_25 sn87_25 11.551961
Rsp86_26 sp86_26 sp87_26 11.551961
Rsn86_26 sn86_26 sn87_26 11.551961
Rsp86_27 sp86_27 sp87_27 11.551961
Rsn86_27 sn86_27 sn87_27 11.551961
Rsp86_28 sp86_28 sp87_28 11.551961
Rsn86_28 sn86_28 sn87_28 11.551961
Rsp86_29 sp86_29 sp87_29 11.551961
Rsn86_29 sn86_29 sn87_29 11.551961
Rsp86_30 sp86_30 sp87_30 11.551961
Rsn86_30 sn86_30 sn87_30 11.551961
Rsp86_31 sp86_31 sp87_31 11.551961
Rsn86_31 sn86_31 sn87_31 11.551961
Rsp86_32 sp86_32 sp87_32 11.551961
Rsn86_32 sn86_32 sn87_32 11.551961
Rsp86_33 sp86_33 sp87_33 11.551961
Rsn86_33 sn86_33 sn87_33 11.551961
Rsp86_34 sp86_34 sp87_34 11.551961
Rsn86_34 sn86_34 sn87_34 11.551961
Rsp86_35 sp86_35 sp87_35 11.551961
Rsn86_35 sn86_35 sn87_35 11.551961
Rsp86_36 sp86_36 sp87_36 11.551961
Rsn86_36 sn86_36 sn87_36 11.551961
Rsp86_37 sp86_37 sp87_37 11.551961
Rsn86_37 sn86_37 sn87_37 11.551961
Rsp86_38 sp86_38 sp87_38 11.551961
Rsn86_38 sn86_38 sn87_38 11.551961
Rsp86_39 sp86_39 sp87_39 11.551961
Rsn86_39 sn86_39 sn87_39 11.551961
Rsp86_40 sp86_40 sp87_40 11.551961
Rsn86_40 sn86_40 sn87_40 11.551961
Rsp86_41 sp86_41 sp87_41 11.551961
Rsn86_41 sn86_41 sn87_41 11.551961
Rsp86_42 sp86_42 sp87_42 11.551961
Rsn86_42 sn86_42 sn87_42 11.551961
Rsp86_43 sp86_43 sp87_43 11.551961
Rsn86_43 sn86_43 sn87_43 11.551961
Rsp86_44 sp86_44 sp87_44 11.551961
Rsn86_44 sn86_44 sn87_44 11.551961
Rsp86_45 sp86_45 sp87_45 11.551961
Rsn86_45 sn86_45 sn87_45 11.551961
Rsp86_46 sp86_46 sp87_46 11.551961
Rsn86_46 sn86_46 sn87_46 11.551961
Rsp86_47 sp86_47 sp87_47 11.551961
Rsn86_47 sn86_47 sn87_47 11.551961
Rsp86_48 sp86_48 sp87_48 11.551961
Rsn86_48 sn86_48 sn87_48 11.551961
Rsp86_49 sp86_49 sp87_49 11.551961
Rsn86_49 sn86_49 sn87_49 11.551961
Rsp86_50 sp86_50 sp87_50 11.551961
Rsn86_50 sn86_50 sn87_50 11.551961
Rsp86_51 sp86_51 sp87_51 11.551961
Rsn86_51 sn86_51 sn87_51 11.551961
Rsp86_52 sp86_52 sp87_52 11.551961
Rsn86_52 sn86_52 sn87_52 11.551961
Rsp86_53 sp86_53 sp87_53 11.551961
Rsn86_53 sn86_53 sn87_53 11.551961
Rsp86_54 sp86_54 sp87_54 11.551961
Rsn86_54 sn86_54 sn87_54 11.551961
Rsp86_55 sp86_55 sp87_55 11.551961
Rsn86_55 sn86_55 sn87_55 11.551961
Rsp86_56 sp86_56 sp87_56 11.551961
Rsn86_56 sn86_56 sn87_56 11.551961
Rsp86_57 sp86_57 sp87_57 11.551961
Rsn86_57 sn86_57 sn87_57 11.551961
Rsp86_58 sp86_58 sp87_58 11.551961
Rsn86_58 sn86_58 sn87_58 11.551961
Rsp86_59 sp86_59 sp87_59 11.551961
Rsn86_59 sn86_59 sn87_59 11.551961
Rsp86_60 sp86_60 sp87_60 11.551961
Rsn86_60 sn86_60 sn87_60 11.551961
Rsp86_61 sp86_61 sp87_61 11.551961
Rsn86_61 sn86_61 sn87_61 11.551961
Rsp86_62 sp86_62 sp87_62 11.551961
Rsn86_62 sn86_62 sn87_62 11.551961
Rsp86_63 sp86_63 sp87_63 11.551961
Rsn86_63 sn86_63 sn87_63 11.551961
Rsp86_64 sp86_64 sp87_64 11.551961
Rsn86_64 sn86_64 sn87_64 11.551961
Rsp86_65 sp86_65 sp87_65 11.551961
Rsn86_65 sn86_65 sn87_65 11.551961
Rsp86_66 sp86_66 sp87_66 11.551961
Rsn86_66 sn86_66 sn87_66 11.551961
Rsp86_67 sp86_67 sp87_67 11.551961
Rsn86_67 sn86_67 sn87_67 11.551961
Rsp86_68 sp86_68 sp87_68 11.551961
Rsn86_68 sn86_68 sn87_68 11.551961
Rsp86_69 sp86_69 sp87_69 11.551961
Rsn86_69 sn86_69 sn87_69 11.551961
Rsp86_70 sp86_70 sp87_70 11.551961
Rsn86_70 sn86_70 sn87_70 11.551961
Rsp86_71 sp86_71 sp87_71 11.551961
Rsn86_71 sn86_71 sn87_71 11.551961
Rsp86_72 sp86_72 sp87_72 11.551961
Rsn86_72 sn86_72 sn87_72 11.551961
Rsp86_73 sp86_73 sp87_73 11.551961
Rsn86_73 sn86_73 sn87_73 11.551961
Rsp86_74 sp86_74 sp87_74 11.551961
Rsn86_74 sn86_74 sn87_74 11.551961
Rsp86_75 sp86_75 sp87_75 11.551961
Rsn86_75 sn86_75 sn87_75 11.551961
Rsp86_76 sp86_76 sp87_76 11.551961
Rsn86_76 sn86_76 sn87_76 11.551961
Rsp86_77 sp86_77 sp87_77 11.551961
Rsn86_77 sn86_77 sn87_77 11.551961
Rsp86_78 sp86_78 sp87_78 11.551961
Rsn86_78 sn86_78 sn87_78 11.551961
Rsp86_79 sp86_79 sp87_79 11.551961
Rsn86_79 sn86_79 sn87_79 11.551961
Rsp86_80 sp86_80 sp87_80 11.551961
Rsn86_80 sn86_80 sn87_80 11.551961
Rsp86_81 sp86_81 sp87_81 11.551961
Rsn86_81 sn86_81 sn87_81 11.551961
Rsp86_82 sp86_82 sp87_82 11.551961
Rsn86_82 sn86_82 sn87_82 11.551961
Rsp86_83 sp86_83 sp87_83 11.551961
Rsn86_83 sn86_83 sn87_83 11.551961
Rsp86_84 sp86_84 sp87_84 11.551961
Rsn86_84 sn86_84 sn87_84 11.551961
Rsp87_1 sp87_1 sp88_1 11.551961
Rsn87_1 sn87_1 sn88_1 11.551961
Rsp87_2 sp87_2 sp88_2 11.551961
Rsn87_2 sn87_2 sn88_2 11.551961
Rsp87_3 sp87_3 sp88_3 11.551961
Rsn87_3 sn87_3 sn88_3 11.551961
Rsp87_4 sp87_4 sp88_4 11.551961
Rsn87_4 sn87_4 sn88_4 11.551961
Rsp87_5 sp87_5 sp88_5 11.551961
Rsn87_5 sn87_5 sn88_5 11.551961
Rsp87_6 sp87_6 sp88_6 11.551961
Rsn87_6 sn87_6 sn88_6 11.551961
Rsp87_7 sp87_7 sp88_7 11.551961
Rsn87_7 sn87_7 sn88_7 11.551961
Rsp87_8 sp87_8 sp88_8 11.551961
Rsn87_8 sn87_8 sn88_8 11.551961
Rsp87_9 sp87_9 sp88_9 11.551961
Rsn87_9 sn87_9 sn88_9 11.551961
Rsp87_10 sp87_10 sp88_10 11.551961
Rsn87_10 sn87_10 sn88_10 11.551961
Rsp87_11 sp87_11 sp88_11 11.551961
Rsn87_11 sn87_11 sn88_11 11.551961
Rsp87_12 sp87_12 sp88_12 11.551961
Rsn87_12 sn87_12 sn88_12 11.551961
Rsp87_13 sp87_13 sp88_13 11.551961
Rsn87_13 sn87_13 sn88_13 11.551961
Rsp87_14 sp87_14 sp88_14 11.551961
Rsn87_14 sn87_14 sn88_14 11.551961
Rsp87_15 sp87_15 sp88_15 11.551961
Rsn87_15 sn87_15 sn88_15 11.551961
Rsp87_16 sp87_16 sp88_16 11.551961
Rsn87_16 sn87_16 sn88_16 11.551961
Rsp87_17 sp87_17 sp88_17 11.551961
Rsn87_17 sn87_17 sn88_17 11.551961
Rsp87_18 sp87_18 sp88_18 11.551961
Rsn87_18 sn87_18 sn88_18 11.551961
Rsp87_19 sp87_19 sp88_19 11.551961
Rsn87_19 sn87_19 sn88_19 11.551961
Rsp87_20 sp87_20 sp88_20 11.551961
Rsn87_20 sn87_20 sn88_20 11.551961
Rsp87_21 sp87_21 sp88_21 11.551961
Rsn87_21 sn87_21 sn88_21 11.551961
Rsp87_22 sp87_22 sp88_22 11.551961
Rsn87_22 sn87_22 sn88_22 11.551961
Rsp87_23 sp87_23 sp88_23 11.551961
Rsn87_23 sn87_23 sn88_23 11.551961
Rsp87_24 sp87_24 sp88_24 11.551961
Rsn87_24 sn87_24 sn88_24 11.551961
Rsp87_25 sp87_25 sp88_25 11.551961
Rsn87_25 sn87_25 sn88_25 11.551961
Rsp87_26 sp87_26 sp88_26 11.551961
Rsn87_26 sn87_26 sn88_26 11.551961
Rsp87_27 sp87_27 sp88_27 11.551961
Rsn87_27 sn87_27 sn88_27 11.551961
Rsp87_28 sp87_28 sp88_28 11.551961
Rsn87_28 sn87_28 sn88_28 11.551961
Rsp87_29 sp87_29 sp88_29 11.551961
Rsn87_29 sn87_29 sn88_29 11.551961
Rsp87_30 sp87_30 sp88_30 11.551961
Rsn87_30 sn87_30 sn88_30 11.551961
Rsp87_31 sp87_31 sp88_31 11.551961
Rsn87_31 sn87_31 sn88_31 11.551961
Rsp87_32 sp87_32 sp88_32 11.551961
Rsn87_32 sn87_32 sn88_32 11.551961
Rsp87_33 sp87_33 sp88_33 11.551961
Rsn87_33 sn87_33 sn88_33 11.551961
Rsp87_34 sp87_34 sp88_34 11.551961
Rsn87_34 sn87_34 sn88_34 11.551961
Rsp87_35 sp87_35 sp88_35 11.551961
Rsn87_35 sn87_35 sn88_35 11.551961
Rsp87_36 sp87_36 sp88_36 11.551961
Rsn87_36 sn87_36 sn88_36 11.551961
Rsp87_37 sp87_37 sp88_37 11.551961
Rsn87_37 sn87_37 sn88_37 11.551961
Rsp87_38 sp87_38 sp88_38 11.551961
Rsn87_38 sn87_38 sn88_38 11.551961
Rsp87_39 sp87_39 sp88_39 11.551961
Rsn87_39 sn87_39 sn88_39 11.551961
Rsp87_40 sp87_40 sp88_40 11.551961
Rsn87_40 sn87_40 sn88_40 11.551961
Rsp87_41 sp87_41 sp88_41 11.551961
Rsn87_41 sn87_41 sn88_41 11.551961
Rsp87_42 sp87_42 sp88_42 11.551961
Rsn87_42 sn87_42 sn88_42 11.551961
Rsp87_43 sp87_43 sp88_43 11.551961
Rsn87_43 sn87_43 sn88_43 11.551961
Rsp87_44 sp87_44 sp88_44 11.551961
Rsn87_44 sn87_44 sn88_44 11.551961
Rsp87_45 sp87_45 sp88_45 11.551961
Rsn87_45 sn87_45 sn88_45 11.551961
Rsp87_46 sp87_46 sp88_46 11.551961
Rsn87_46 sn87_46 sn88_46 11.551961
Rsp87_47 sp87_47 sp88_47 11.551961
Rsn87_47 sn87_47 sn88_47 11.551961
Rsp87_48 sp87_48 sp88_48 11.551961
Rsn87_48 sn87_48 sn88_48 11.551961
Rsp87_49 sp87_49 sp88_49 11.551961
Rsn87_49 sn87_49 sn88_49 11.551961
Rsp87_50 sp87_50 sp88_50 11.551961
Rsn87_50 sn87_50 sn88_50 11.551961
Rsp87_51 sp87_51 sp88_51 11.551961
Rsn87_51 sn87_51 sn88_51 11.551961
Rsp87_52 sp87_52 sp88_52 11.551961
Rsn87_52 sn87_52 sn88_52 11.551961
Rsp87_53 sp87_53 sp88_53 11.551961
Rsn87_53 sn87_53 sn88_53 11.551961
Rsp87_54 sp87_54 sp88_54 11.551961
Rsn87_54 sn87_54 sn88_54 11.551961
Rsp87_55 sp87_55 sp88_55 11.551961
Rsn87_55 sn87_55 sn88_55 11.551961
Rsp87_56 sp87_56 sp88_56 11.551961
Rsn87_56 sn87_56 sn88_56 11.551961
Rsp87_57 sp87_57 sp88_57 11.551961
Rsn87_57 sn87_57 sn88_57 11.551961
Rsp87_58 sp87_58 sp88_58 11.551961
Rsn87_58 sn87_58 sn88_58 11.551961
Rsp87_59 sp87_59 sp88_59 11.551961
Rsn87_59 sn87_59 sn88_59 11.551961
Rsp87_60 sp87_60 sp88_60 11.551961
Rsn87_60 sn87_60 sn88_60 11.551961
Rsp87_61 sp87_61 sp88_61 11.551961
Rsn87_61 sn87_61 sn88_61 11.551961
Rsp87_62 sp87_62 sp88_62 11.551961
Rsn87_62 sn87_62 sn88_62 11.551961
Rsp87_63 sp87_63 sp88_63 11.551961
Rsn87_63 sn87_63 sn88_63 11.551961
Rsp87_64 sp87_64 sp88_64 11.551961
Rsn87_64 sn87_64 sn88_64 11.551961
Rsp87_65 sp87_65 sp88_65 11.551961
Rsn87_65 sn87_65 sn88_65 11.551961
Rsp87_66 sp87_66 sp88_66 11.551961
Rsn87_66 sn87_66 sn88_66 11.551961
Rsp87_67 sp87_67 sp88_67 11.551961
Rsn87_67 sn87_67 sn88_67 11.551961
Rsp87_68 sp87_68 sp88_68 11.551961
Rsn87_68 sn87_68 sn88_68 11.551961
Rsp87_69 sp87_69 sp88_69 11.551961
Rsn87_69 sn87_69 sn88_69 11.551961
Rsp87_70 sp87_70 sp88_70 11.551961
Rsn87_70 sn87_70 sn88_70 11.551961
Rsp87_71 sp87_71 sp88_71 11.551961
Rsn87_71 sn87_71 sn88_71 11.551961
Rsp87_72 sp87_72 sp88_72 11.551961
Rsn87_72 sn87_72 sn88_72 11.551961
Rsp87_73 sp87_73 sp88_73 11.551961
Rsn87_73 sn87_73 sn88_73 11.551961
Rsp87_74 sp87_74 sp88_74 11.551961
Rsn87_74 sn87_74 sn88_74 11.551961
Rsp87_75 sp87_75 sp88_75 11.551961
Rsn87_75 sn87_75 sn88_75 11.551961
Rsp87_76 sp87_76 sp88_76 11.551961
Rsn87_76 sn87_76 sn88_76 11.551961
Rsp87_77 sp87_77 sp88_77 11.551961
Rsn87_77 sn87_77 sn88_77 11.551961
Rsp87_78 sp87_78 sp88_78 11.551961
Rsn87_78 sn87_78 sn88_78 11.551961
Rsp87_79 sp87_79 sp88_79 11.551961
Rsn87_79 sn87_79 sn88_79 11.551961
Rsp87_80 sp87_80 sp88_80 11.551961
Rsn87_80 sn87_80 sn88_80 11.551961
Rsp87_81 sp87_81 sp88_81 11.551961
Rsn87_81 sn87_81 sn88_81 11.551961
Rsp87_82 sp87_82 sp88_82 11.551961
Rsn87_82 sn87_82 sn88_82 11.551961
Rsp87_83 sp87_83 sp88_83 11.551961
Rsn87_83 sn87_83 sn88_83 11.551961
Rsp87_84 sp87_84 sp88_84 11.551961
Rsn87_84 sn87_84 sn88_84 11.551961
Rsp88_1 sp88_1 sp89_1 11.551961
Rsn88_1 sn88_1 sn89_1 11.551961
Rsp88_2 sp88_2 sp89_2 11.551961
Rsn88_2 sn88_2 sn89_2 11.551961
Rsp88_3 sp88_3 sp89_3 11.551961
Rsn88_3 sn88_3 sn89_3 11.551961
Rsp88_4 sp88_4 sp89_4 11.551961
Rsn88_4 sn88_4 sn89_4 11.551961
Rsp88_5 sp88_5 sp89_5 11.551961
Rsn88_5 sn88_5 sn89_5 11.551961
Rsp88_6 sp88_6 sp89_6 11.551961
Rsn88_6 sn88_6 sn89_6 11.551961
Rsp88_7 sp88_7 sp89_7 11.551961
Rsn88_7 sn88_7 sn89_7 11.551961
Rsp88_8 sp88_8 sp89_8 11.551961
Rsn88_8 sn88_8 sn89_8 11.551961
Rsp88_9 sp88_9 sp89_9 11.551961
Rsn88_9 sn88_9 sn89_9 11.551961
Rsp88_10 sp88_10 sp89_10 11.551961
Rsn88_10 sn88_10 sn89_10 11.551961
Rsp88_11 sp88_11 sp89_11 11.551961
Rsn88_11 sn88_11 sn89_11 11.551961
Rsp88_12 sp88_12 sp89_12 11.551961
Rsn88_12 sn88_12 sn89_12 11.551961
Rsp88_13 sp88_13 sp89_13 11.551961
Rsn88_13 sn88_13 sn89_13 11.551961
Rsp88_14 sp88_14 sp89_14 11.551961
Rsn88_14 sn88_14 sn89_14 11.551961
Rsp88_15 sp88_15 sp89_15 11.551961
Rsn88_15 sn88_15 sn89_15 11.551961
Rsp88_16 sp88_16 sp89_16 11.551961
Rsn88_16 sn88_16 sn89_16 11.551961
Rsp88_17 sp88_17 sp89_17 11.551961
Rsn88_17 sn88_17 sn89_17 11.551961
Rsp88_18 sp88_18 sp89_18 11.551961
Rsn88_18 sn88_18 sn89_18 11.551961
Rsp88_19 sp88_19 sp89_19 11.551961
Rsn88_19 sn88_19 sn89_19 11.551961
Rsp88_20 sp88_20 sp89_20 11.551961
Rsn88_20 sn88_20 sn89_20 11.551961
Rsp88_21 sp88_21 sp89_21 11.551961
Rsn88_21 sn88_21 sn89_21 11.551961
Rsp88_22 sp88_22 sp89_22 11.551961
Rsn88_22 sn88_22 sn89_22 11.551961
Rsp88_23 sp88_23 sp89_23 11.551961
Rsn88_23 sn88_23 sn89_23 11.551961
Rsp88_24 sp88_24 sp89_24 11.551961
Rsn88_24 sn88_24 sn89_24 11.551961
Rsp88_25 sp88_25 sp89_25 11.551961
Rsn88_25 sn88_25 sn89_25 11.551961
Rsp88_26 sp88_26 sp89_26 11.551961
Rsn88_26 sn88_26 sn89_26 11.551961
Rsp88_27 sp88_27 sp89_27 11.551961
Rsn88_27 sn88_27 sn89_27 11.551961
Rsp88_28 sp88_28 sp89_28 11.551961
Rsn88_28 sn88_28 sn89_28 11.551961
Rsp88_29 sp88_29 sp89_29 11.551961
Rsn88_29 sn88_29 sn89_29 11.551961
Rsp88_30 sp88_30 sp89_30 11.551961
Rsn88_30 sn88_30 sn89_30 11.551961
Rsp88_31 sp88_31 sp89_31 11.551961
Rsn88_31 sn88_31 sn89_31 11.551961
Rsp88_32 sp88_32 sp89_32 11.551961
Rsn88_32 sn88_32 sn89_32 11.551961
Rsp88_33 sp88_33 sp89_33 11.551961
Rsn88_33 sn88_33 sn89_33 11.551961
Rsp88_34 sp88_34 sp89_34 11.551961
Rsn88_34 sn88_34 sn89_34 11.551961
Rsp88_35 sp88_35 sp89_35 11.551961
Rsn88_35 sn88_35 sn89_35 11.551961
Rsp88_36 sp88_36 sp89_36 11.551961
Rsn88_36 sn88_36 sn89_36 11.551961
Rsp88_37 sp88_37 sp89_37 11.551961
Rsn88_37 sn88_37 sn89_37 11.551961
Rsp88_38 sp88_38 sp89_38 11.551961
Rsn88_38 sn88_38 sn89_38 11.551961
Rsp88_39 sp88_39 sp89_39 11.551961
Rsn88_39 sn88_39 sn89_39 11.551961
Rsp88_40 sp88_40 sp89_40 11.551961
Rsn88_40 sn88_40 sn89_40 11.551961
Rsp88_41 sp88_41 sp89_41 11.551961
Rsn88_41 sn88_41 sn89_41 11.551961
Rsp88_42 sp88_42 sp89_42 11.551961
Rsn88_42 sn88_42 sn89_42 11.551961
Rsp88_43 sp88_43 sp89_43 11.551961
Rsn88_43 sn88_43 sn89_43 11.551961
Rsp88_44 sp88_44 sp89_44 11.551961
Rsn88_44 sn88_44 sn89_44 11.551961
Rsp88_45 sp88_45 sp89_45 11.551961
Rsn88_45 sn88_45 sn89_45 11.551961
Rsp88_46 sp88_46 sp89_46 11.551961
Rsn88_46 sn88_46 sn89_46 11.551961
Rsp88_47 sp88_47 sp89_47 11.551961
Rsn88_47 sn88_47 sn89_47 11.551961
Rsp88_48 sp88_48 sp89_48 11.551961
Rsn88_48 sn88_48 sn89_48 11.551961
Rsp88_49 sp88_49 sp89_49 11.551961
Rsn88_49 sn88_49 sn89_49 11.551961
Rsp88_50 sp88_50 sp89_50 11.551961
Rsn88_50 sn88_50 sn89_50 11.551961
Rsp88_51 sp88_51 sp89_51 11.551961
Rsn88_51 sn88_51 sn89_51 11.551961
Rsp88_52 sp88_52 sp89_52 11.551961
Rsn88_52 sn88_52 sn89_52 11.551961
Rsp88_53 sp88_53 sp89_53 11.551961
Rsn88_53 sn88_53 sn89_53 11.551961
Rsp88_54 sp88_54 sp89_54 11.551961
Rsn88_54 sn88_54 sn89_54 11.551961
Rsp88_55 sp88_55 sp89_55 11.551961
Rsn88_55 sn88_55 sn89_55 11.551961
Rsp88_56 sp88_56 sp89_56 11.551961
Rsn88_56 sn88_56 sn89_56 11.551961
Rsp88_57 sp88_57 sp89_57 11.551961
Rsn88_57 sn88_57 sn89_57 11.551961
Rsp88_58 sp88_58 sp89_58 11.551961
Rsn88_58 sn88_58 sn89_58 11.551961
Rsp88_59 sp88_59 sp89_59 11.551961
Rsn88_59 sn88_59 sn89_59 11.551961
Rsp88_60 sp88_60 sp89_60 11.551961
Rsn88_60 sn88_60 sn89_60 11.551961
Rsp88_61 sp88_61 sp89_61 11.551961
Rsn88_61 sn88_61 sn89_61 11.551961
Rsp88_62 sp88_62 sp89_62 11.551961
Rsn88_62 sn88_62 sn89_62 11.551961
Rsp88_63 sp88_63 sp89_63 11.551961
Rsn88_63 sn88_63 sn89_63 11.551961
Rsp88_64 sp88_64 sp89_64 11.551961
Rsn88_64 sn88_64 sn89_64 11.551961
Rsp88_65 sp88_65 sp89_65 11.551961
Rsn88_65 sn88_65 sn89_65 11.551961
Rsp88_66 sp88_66 sp89_66 11.551961
Rsn88_66 sn88_66 sn89_66 11.551961
Rsp88_67 sp88_67 sp89_67 11.551961
Rsn88_67 sn88_67 sn89_67 11.551961
Rsp88_68 sp88_68 sp89_68 11.551961
Rsn88_68 sn88_68 sn89_68 11.551961
Rsp88_69 sp88_69 sp89_69 11.551961
Rsn88_69 sn88_69 sn89_69 11.551961
Rsp88_70 sp88_70 sp89_70 11.551961
Rsn88_70 sn88_70 sn89_70 11.551961
Rsp88_71 sp88_71 sp89_71 11.551961
Rsn88_71 sn88_71 sn89_71 11.551961
Rsp88_72 sp88_72 sp89_72 11.551961
Rsn88_72 sn88_72 sn89_72 11.551961
Rsp88_73 sp88_73 sp89_73 11.551961
Rsn88_73 sn88_73 sn89_73 11.551961
Rsp88_74 sp88_74 sp89_74 11.551961
Rsn88_74 sn88_74 sn89_74 11.551961
Rsp88_75 sp88_75 sp89_75 11.551961
Rsn88_75 sn88_75 sn89_75 11.551961
Rsp88_76 sp88_76 sp89_76 11.551961
Rsn88_76 sn88_76 sn89_76 11.551961
Rsp88_77 sp88_77 sp89_77 11.551961
Rsn88_77 sn88_77 sn89_77 11.551961
Rsp88_78 sp88_78 sp89_78 11.551961
Rsn88_78 sn88_78 sn89_78 11.551961
Rsp88_79 sp88_79 sp89_79 11.551961
Rsn88_79 sn88_79 sn89_79 11.551961
Rsp88_80 sp88_80 sp89_80 11.551961
Rsn88_80 sn88_80 sn89_80 11.551961
Rsp88_81 sp88_81 sp89_81 11.551961
Rsn88_81 sn88_81 sn89_81 11.551961
Rsp88_82 sp88_82 sp89_82 11.551961
Rsn88_82 sn88_82 sn89_82 11.551961
Rsp88_83 sp88_83 sp89_83 11.551961
Rsn88_83 sn88_83 sn89_83 11.551961
Rsp88_84 sp88_84 sp89_84 11.551961
Rsn88_84 sn88_84 sn89_84 11.551961
Rsp89_1 sp89_1 sp90_1 11.551961
Rsn89_1 sn89_1 sn90_1 11.551961
Rsp89_2 sp89_2 sp90_2 11.551961
Rsn89_2 sn89_2 sn90_2 11.551961
Rsp89_3 sp89_3 sp90_3 11.551961
Rsn89_3 sn89_3 sn90_3 11.551961
Rsp89_4 sp89_4 sp90_4 11.551961
Rsn89_4 sn89_4 sn90_4 11.551961
Rsp89_5 sp89_5 sp90_5 11.551961
Rsn89_5 sn89_5 sn90_5 11.551961
Rsp89_6 sp89_6 sp90_6 11.551961
Rsn89_6 sn89_6 sn90_6 11.551961
Rsp89_7 sp89_7 sp90_7 11.551961
Rsn89_7 sn89_7 sn90_7 11.551961
Rsp89_8 sp89_8 sp90_8 11.551961
Rsn89_8 sn89_8 sn90_8 11.551961
Rsp89_9 sp89_9 sp90_9 11.551961
Rsn89_9 sn89_9 sn90_9 11.551961
Rsp89_10 sp89_10 sp90_10 11.551961
Rsn89_10 sn89_10 sn90_10 11.551961
Rsp89_11 sp89_11 sp90_11 11.551961
Rsn89_11 sn89_11 sn90_11 11.551961
Rsp89_12 sp89_12 sp90_12 11.551961
Rsn89_12 sn89_12 sn90_12 11.551961
Rsp89_13 sp89_13 sp90_13 11.551961
Rsn89_13 sn89_13 sn90_13 11.551961
Rsp89_14 sp89_14 sp90_14 11.551961
Rsn89_14 sn89_14 sn90_14 11.551961
Rsp89_15 sp89_15 sp90_15 11.551961
Rsn89_15 sn89_15 sn90_15 11.551961
Rsp89_16 sp89_16 sp90_16 11.551961
Rsn89_16 sn89_16 sn90_16 11.551961
Rsp89_17 sp89_17 sp90_17 11.551961
Rsn89_17 sn89_17 sn90_17 11.551961
Rsp89_18 sp89_18 sp90_18 11.551961
Rsn89_18 sn89_18 sn90_18 11.551961
Rsp89_19 sp89_19 sp90_19 11.551961
Rsn89_19 sn89_19 sn90_19 11.551961
Rsp89_20 sp89_20 sp90_20 11.551961
Rsn89_20 sn89_20 sn90_20 11.551961
Rsp89_21 sp89_21 sp90_21 11.551961
Rsn89_21 sn89_21 sn90_21 11.551961
Rsp89_22 sp89_22 sp90_22 11.551961
Rsn89_22 sn89_22 sn90_22 11.551961
Rsp89_23 sp89_23 sp90_23 11.551961
Rsn89_23 sn89_23 sn90_23 11.551961
Rsp89_24 sp89_24 sp90_24 11.551961
Rsn89_24 sn89_24 sn90_24 11.551961
Rsp89_25 sp89_25 sp90_25 11.551961
Rsn89_25 sn89_25 sn90_25 11.551961
Rsp89_26 sp89_26 sp90_26 11.551961
Rsn89_26 sn89_26 sn90_26 11.551961
Rsp89_27 sp89_27 sp90_27 11.551961
Rsn89_27 sn89_27 sn90_27 11.551961
Rsp89_28 sp89_28 sp90_28 11.551961
Rsn89_28 sn89_28 sn90_28 11.551961
Rsp89_29 sp89_29 sp90_29 11.551961
Rsn89_29 sn89_29 sn90_29 11.551961
Rsp89_30 sp89_30 sp90_30 11.551961
Rsn89_30 sn89_30 sn90_30 11.551961
Rsp89_31 sp89_31 sp90_31 11.551961
Rsn89_31 sn89_31 sn90_31 11.551961
Rsp89_32 sp89_32 sp90_32 11.551961
Rsn89_32 sn89_32 sn90_32 11.551961
Rsp89_33 sp89_33 sp90_33 11.551961
Rsn89_33 sn89_33 sn90_33 11.551961
Rsp89_34 sp89_34 sp90_34 11.551961
Rsn89_34 sn89_34 sn90_34 11.551961
Rsp89_35 sp89_35 sp90_35 11.551961
Rsn89_35 sn89_35 sn90_35 11.551961
Rsp89_36 sp89_36 sp90_36 11.551961
Rsn89_36 sn89_36 sn90_36 11.551961
Rsp89_37 sp89_37 sp90_37 11.551961
Rsn89_37 sn89_37 sn90_37 11.551961
Rsp89_38 sp89_38 sp90_38 11.551961
Rsn89_38 sn89_38 sn90_38 11.551961
Rsp89_39 sp89_39 sp90_39 11.551961
Rsn89_39 sn89_39 sn90_39 11.551961
Rsp89_40 sp89_40 sp90_40 11.551961
Rsn89_40 sn89_40 sn90_40 11.551961
Rsp89_41 sp89_41 sp90_41 11.551961
Rsn89_41 sn89_41 sn90_41 11.551961
Rsp89_42 sp89_42 sp90_42 11.551961
Rsn89_42 sn89_42 sn90_42 11.551961
Rsp89_43 sp89_43 sp90_43 11.551961
Rsn89_43 sn89_43 sn90_43 11.551961
Rsp89_44 sp89_44 sp90_44 11.551961
Rsn89_44 sn89_44 sn90_44 11.551961
Rsp89_45 sp89_45 sp90_45 11.551961
Rsn89_45 sn89_45 sn90_45 11.551961
Rsp89_46 sp89_46 sp90_46 11.551961
Rsn89_46 sn89_46 sn90_46 11.551961
Rsp89_47 sp89_47 sp90_47 11.551961
Rsn89_47 sn89_47 sn90_47 11.551961
Rsp89_48 sp89_48 sp90_48 11.551961
Rsn89_48 sn89_48 sn90_48 11.551961
Rsp89_49 sp89_49 sp90_49 11.551961
Rsn89_49 sn89_49 sn90_49 11.551961
Rsp89_50 sp89_50 sp90_50 11.551961
Rsn89_50 sn89_50 sn90_50 11.551961
Rsp89_51 sp89_51 sp90_51 11.551961
Rsn89_51 sn89_51 sn90_51 11.551961
Rsp89_52 sp89_52 sp90_52 11.551961
Rsn89_52 sn89_52 sn90_52 11.551961
Rsp89_53 sp89_53 sp90_53 11.551961
Rsn89_53 sn89_53 sn90_53 11.551961
Rsp89_54 sp89_54 sp90_54 11.551961
Rsn89_54 sn89_54 sn90_54 11.551961
Rsp89_55 sp89_55 sp90_55 11.551961
Rsn89_55 sn89_55 sn90_55 11.551961
Rsp89_56 sp89_56 sp90_56 11.551961
Rsn89_56 sn89_56 sn90_56 11.551961
Rsp89_57 sp89_57 sp90_57 11.551961
Rsn89_57 sn89_57 sn90_57 11.551961
Rsp89_58 sp89_58 sp90_58 11.551961
Rsn89_58 sn89_58 sn90_58 11.551961
Rsp89_59 sp89_59 sp90_59 11.551961
Rsn89_59 sn89_59 sn90_59 11.551961
Rsp89_60 sp89_60 sp90_60 11.551961
Rsn89_60 sn89_60 sn90_60 11.551961
Rsp89_61 sp89_61 sp90_61 11.551961
Rsn89_61 sn89_61 sn90_61 11.551961
Rsp89_62 sp89_62 sp90_62 11.551961
Rsn89_62 sn89_62 sn90_62 11.551961
Rsp89_63 sp89_63 sp90_63 11.551961
Rsn89_63 sn89_63 sn90_63 11.551961
Rsp89_64 sp89_64 sp90_64 11.551961
Rsn89_64 sn89_64 sn90_64 11.551961
Rsp89_65 sp89_65 sp90_65 11.551961
Rsn89_65 sn89_65 sn90_65 11.551961
Rsp89_66 sp89_66 sp90_66 11.551961
Rsn89_66 sn89_66 sn90_66 11.551961
Rsp89_67 sp89_67 sp90_67 11.551961
Rsn89_67 sn89_67 sn90_67 11.551961
Rsp89_68 sp89_68 sp90_68 11.551961
Rsn89_68 sn89_68 sn90_68 11.551961
Rsp89_69 sp89_69 sp90_69 11.551961
Rsn89_69 sn89_69 sn90_69 11.551961
Rsp89_70 sp89_70 sp90_70 11.551961
Rsn89_70 sn89_70 sn90_70 11.551961
Rsp89_71 sp89_71 sp90_71 11.551961
Rsn89_71 sn89_71 sn90_71 11.551961
Rsp89_72 sp89_72 sp90_72 11.551961
Rsn89_72 sn89_72 sn90_72 11.551961
Rsp89_73 sp89_73 sp90_73 11.551961
Rsn89_73 sn89_73 sn90_73 11.551961
Rsp89_74 sp89_74 sp90_74 11.551961
Rsn89_74 sn89_74 sn90_74 11.551961
Rsp89_75 sp89_75 sp90_75 11.551961
Rsn89_75 sn89_75 sn90_75 11.551961
Rsp89_76 sp89_76 sp90_76 11.551961
Rsn89_76 sn89_76 sn90_76 11.551961
Rsp89_77 sp89_77 sp90_77 11.551961
Rsn89_77 sn89_77 sn90_77 11.551961
Rsp89_78 sp89_78 sp90_78 11.551961
Rsn89_78 sn89_78 sn90_78 11.551961
Rsp89_79 sp89_79 sp90_79 11.551961
Rsn89_79 sn89_79 sn90_79 11.551961
Rsp89_80 sp89_80 sp90_80 11.551961
Rsn89_80 sn89_80 sn90_80 11.551961
Rsp89_81 sp89_81 sp90_81 11.551961
Rsn89_81 sn89_81 sn90_81 11.551961
Rsp89_82 sp89_82 sp90_82 11.551961
Rsn89_82 sn89_82 sn90_82 11.551961
Rsp89_83 sp89_83 sp90_83 11.551961
Rsn89_83 sn89_83 sn90_83 11.551961
Rsp89_84 sp89_84 sp90_84 11.551961
Rsn89_84 sn89_84 sn90_84 11.551961
Rsp90_1 sp90_1 sp91_1 11.551961
Rsn90_1 sn90_1 sn91_1 11.551961
Rsp90_2 sp90_2 sp91_2 11.551961
Rsn90_2 sn90_2 sn91_2 11.551961
Rsp90_3 sp90_3 sp91_3 11.551961
Rsn90_3 sn90_3 sn91_3 11.551961
Rsp90_4 sp90_4 sp91_4 11.551961
Rsn90_4 sn90_4 sn91_4 11.551961
Rsp90_5 sp90_5 sp91_5 11.551961
Rsn90_5 sn90_5 sn91_5 11.551961
Rsp90_6 sp90_6 sp91_6 11.551961
Rsn90_6 sn90_6 sn91_6 11.551961
Rsp90_7 sp90_7 sp91_7 11.551961
Rsn90_7 sn90_7 sn91_7 11.551961
Rsp90_8 sp90_8 sp91_8 11.551961
Rsn90_8 sn90_8 sn91_8 11.551961
Rsp90_9 sp90_9 sp91_9 11.551961
Rsn90_9 sn90_9 sn91_9 11.551961
Rsp90_10 sp90_10 sp91_10 11.551961
Rsn90_10 sn90_10 sn91_10 11.551961
Rsp90_11 sp90_11 sp91_11 11.551961
Rsn90_11 sn90_11 sn91_11 11.551961
Rsp90_12 sp90_12 sp91_12 11.551961
Rsn90_12 sn90_12 sn91_12 11.551961
Rsp90_13 sp90_13 sp91_13 11.551961
Rsn90_13 sn90_13 sn91_13 11.551961
Rsp90_14 sp90_14 sp91_14 11.551961
Rsn90_14 sn90_14 sn91_14 11.551961
Rsp90_15 sp90_15 sp91_15 11.551961
Rsn90_15 sn90_15 sn91_15 11.551961
Rsp90_16 sp90_16 sp91_16 11.551961
Rsn90_16 sn90_16 sn91_16 11.551961
Rsp90_17 sp90_17 sp91_17 11.551961
Rsn90_17 sn90_17 sn91_17 11.551961
Rsp90_18 sp90_18 sp91_18 11.551961
Rsn90_18 sn90_18 sn91_18 11.551961
Rsp90_19 sp90_19 sp91_19 11.551961
Rsn90_19 sn90_19 sn91_19 11.551961
Rsp90_20 sp90_20 sp91_20 11.551961
Rsn90_20 sn90_20 sn91_20 11.551961
Rsp90_21 sp90_21 sp91_21 11.551961
Rsn90_21 sn90_21 sn91_21 11.551961
Rsp90_22 sp90_22 sp91_22 11.551961
Rsn90_22 sn90_22 sn91_22 11.551961
Rsp90_23 sp90_23 sp91_23 11.551961
Rsn90_23 sn90_23 sn91_23 11.551961
Rsp90_24 sp90_24 sp91_24 11.551961
Rsn90_24 sn90_24 sn91_24 11.551961
Rsp90_25 sp90_25 sp91_25 11.551961
Rsn90_25 sn90_25 sn91_25 11.551961
Rsp90_26 sp90_26 sp91_26 11.551961
Rsn90_26 sn90_26 sn91_26 11.551961
Rsp90_27 sp90_27 sp91_27 11.551961
Rsn90_27 sn90_27 sn91_27 11.551961
Rsp90_28 sp90_28 sp91_28 11.551961
Rsn90_28 sn90_28 sn91_28 11.551961
Rsp90_29 sp90_29 sp91_29 11.551961
Rsn90_29 sn90_29 sn91_29 11.551961
Rsp90_30 sp90_30 sp91_30 11.551961
Rsn90_30 sn90_30 sn91_30 11.551961
Rsp90_31 sp90_31 sp91_31 11.551961
Rsn90_31 sn90_31 sn91_31 11.551961
Rsp90_32 sp90_32 sp91_32 11.551961
Rsn90_32 sn90_32 sn91_32 11.551961
Rsp90_33 sp90_33 sp91_33 11.551961
Rsn90_33 sn90_33 sn91_33 11.551961
Rsp90_34 sp90_34 sp91_34 11.551961
Rsn90_34 sn90_34 sn91_34 11.551961
Rsp90_35 sp90_35 sp91_35 11.551961
Rsn90_35 sn90_35 sn91_35 11.551961
Rsp90_36 sp90_36 sp91_36 11.551961
Rsn90_36 sn90_36 sn91_36 11.551961
Rsp90_37 sp90_37 sp91_37 11.551961
Rsn90_37 sn90_37 sn91_37 11.551961
Rsp90_38 sp90_38 sp91_38 11.551961
Rsn90_38 sn90_38 sn91_38 11.551961
Rsp90_39 sp90_39 sp91_39 11.551961
Rsn90_39 sn90_39 sn91_39 11.551961
Rsp90_40 sp90_40 sp91_40 11.551961
Rsn90_40 sn90_40 sn91_40 11.551961
Rsp90_41 sp90_41 sp91_41 11.551961
Rsn90_41 sn90_41 sn91_41 11.551961
Rsp90_42 sp90_42 sp91_42 11.551961
Rsn90_42 sn90_42 sn91_42 11.551961
Rsp90_43 sp90_43 sp91_43 11.551961
Rsn90_43 sn90_43 sn91_43 11.551961
Rsp90_44 sp90_44 sp91_44 11.551961
Rsn90_44 sn90_44 sn91_44 11.551961
Rsp90_45 sp90_45 sp91_45 11.551961
Rsn90_45 sn90_45 sn91_45 11.551961
Rsp90_46 sp90_46 sp91_46 11.551961
Rsn90_46 sn90_46 sn91_46 11.551961
Rsp90_47 sp90_47 sp91_47 11.551961
Rsn90_47 sn90_47 sn91_47 11.551961
Rsp90_48 sp90_48 sp91_48 11.551961
Rsn90_48 sn90_48 sn91_48 11.551961
Rsp90_49 sp90_49 sp91_49 11.551961
Rsn90_49 sn90_49 sn91_49 11.551961
Rsp90_50 sp90_50 sp91_50 11.551961
Rsn90_50 sn90_50 sn91_50 11.551961
Rsp90_51 sp90_51 sp91_51 11.551961
Rsn90_51 sn90_51 sn91_51 11.551961
Rsp90_52 sp90_52 sp91_52 11.551961
Rsn90_52 sn90_52 sn91_52 11.551961
Rsp90_53 sp90_53 sp91_53 11.551961
Rsn90_53 sn90_53 sn91_53 11.551961
Rsp90_54 sp90_54 sp91_54 11.551961
Rsn90_54 sn90_54 sn91_54 11.551961
Rsp90_55 sp90_55 sp91_55 11.551961
Rsn90_55 sn90_55 sn91_55 11.551961
Rsp90_56 sp90_56 sp91_56 11.551961
Rsn90_56 sn90_56 sn91_56 11.551961
Rsp90_57 sp90_57 sp91_57 11.551961
Rsn90_57 sn90_57 sn91_57 11.551961
Rsp90_58 sp90_58 sp91_58 11.551961
Rsn90_58 sn90_58 sn91_58 11.551961
Rsp90_59 sp90_59 sp91_59 11.551961
Rsn90_59 sn90_59 sn91_59 11.551961
Rsp90_60 sp90_60 sp91_60 11.551961
Rsn90_60 sn90_60 sn91_60 11.551961
Rsp90_61 sp90_61 sp91_61 11.551961
Rsn90_61 sn90_61 sn91_61 11.551961
Rsp90_62 sp90_62 sp91_62 11.551961
Rsn90_62 sn90_62 sn91_62 11.551961
Rsp90_63 sp90_63 sp91_63 11.551961
Rsn90_63 sn90_63 sn91_63 11.551961
Rsp90_64 sp90_64 sp91_64 11.551961
Rsn90_64 sn90_64 sn91_64 11.551961
Rsp90_65 sp90_65 sp91_65 11.551961
Rsn90_65 sn90_65 sn91_65 11.551961
Rsp90_66 sp90_66 sp91_66 11.551961
Rsn90_66 sn90_66 sn91_66 11.551961
Rsp90_67 sp90_67 sp91_67 11.551961
Rsn90_67 sn90_67 sn91_67 11.551961
Rsp90_68 sp90_68 sp91_68 11.551961
Rsn90_68 sn90_68 sn91_68 11.551961
Rsp90_69 sp90_69 sp91_69 11.551961
Rsn90_69 sn90_69 sn91_69 11.551961
Rsp90_70 sp90_70 sp91_70 11.551961
Rsn90_70 sn90_70 sn91_70 11.551961
Rsp90_71 sp90_71 sp91_71 11.551961
Rsn90_71 sn90_71 sn91_71 11.551961
Rsp90_72 sp90_72 sp91_72 11.551961
Rsn90_72 sn90_72 sn91_72 11.551961
Rsp90_73 sp90_73 sp91_73 11.551961
Rsn90_73 sn90_73 sn91_73 11.551961
Rsp90_74 sp90_74 sp91_74 11.551961
Rsn90_74 sn90_74 sn91_74 11.551961
Rsp90_75 sp90_75 sp91_75 11.551961
Rsn90_75 sn90_75 sn91_75 11.551961
Rsp90_76 sp90_76 sp91_76 11.551961
Rsn90_76 sn90_76 sn91_76 11.551961
Rsp90_77 sp90_77 sp91_77 11.551961
Rsn90_77 sn90_77 sn91_77 11.551961
Rsp90_78 sp90_78 sp91_78 11.551961
Rsn90_78 sn90_78 sn91_78 11.551961
Rsp90_79 sp90_79 sp91_79 11.551961
Rsn90_79 sn90_79 sn91_79 11.551961
Rsp90_80 sp90_80 sp91_80 11.551961
Rsn90_80 sn90_80 sn91_80 11.551961
Rsp90_81 sp90_81 sp91_81 11.551961
Rsn90_81 sn90_81 sn91_81 11.551961
Rsp90_82 sp90_82 sp91_82 11.551961
Rsn90_82 sn90_82 sn91_82 11.551961
Rsp90_83 sp90_83 sp91_83 11.551961
Rsn90_83 sn90_83 sn91_83 11.551961
Rsp90_84 sp90_84 sp91_84 11.551961
Rsn90_84 sn90_84 sn91_84 11.551961
Rsp91_1 sp91_1 sp1_p3 11.551961
Rsn91_1 sn91_1 sn1_p3 11.551961
Rsp91_2 sp91_2 sp2_p3 11.551961
Rsn91_2 sn91_2 sn2_p3 11.551961
Rsp91_3 sp91_3 sp3_p3 11.551961
Rsn91_3 sn91_3 sn3_p3 11.551961
Rsp91_4 sp91_4 sp4_p3 11.551961
Rsn91_4 sn91_4 sn4_p3 11.551961
Rsp91_5 sp91_5 sp5_p3 11.551961
Rsn91_5 sn91_5 sn5_p3 11.551961
Rsp91_6 sp91_6 sp6_p3 11.551961
Rsn91_6 sn91_6 sn6_p3 11.551961
Rsp91_7 sp91_7 sp7_p3 11.551961
Rsn91_7 sn91_7 sn7_p3 11.551961
Rsp91_8 sp91_8 sp8_p3 11.551961
Rsn91_8 sn91_8 sn8_p3 11.551961
Rsp91_9 sp91_9 sp9_p3 11.551961
Rsn91_9 sn91_9 sn9_p3 11.551961
Rsp91_10 sp91_10 sp10_p3 11.551961
Rsn91_10 sn91_10 sn10_p3 11.551961
Rsp91_11 sp91_11 sp11_p3 11.551961
Rsn91_11 sn91_11 sn11_p3 11.551961
Rsp91_12 sp91_12 sp12_p3 11.551961
Rsn91_12 sn91_12 sn12_p3 11.551961
Rsp91_13 sp91_13 sp13_p3 11.551961
Rsn91_13 sn91_13 sn13_p3 11.551961
Rsp91_14 sp91_14 sp14_p3 11.551961
Rsn91_14 sn91_14 sn14_p3 11.551961
Rsp91_15 sp91_15 sp15_p3 11.551961
Rsn91_15 sn91_15 sn15_p3 11.551961
Rsp91_16 sp91_16 sp16_p3 11.551961
Rsn91_16 sn91_16 sn16_p3 11.551961
Rsp91_17 sp91_17 sp17_p3 11.551961
Rsn91_17 sn91_17 sn17_p3 11.551961
Rsp91_18 sp91_18 sp18_p3 11.551961
Rsn91_18 sn91_18 sn18_p3 11.551961
Rsp91_19 sp91_19 sp19_p3 11.551961
Rsn91_19 sn91_19 sn19_p3 11.551961
Rsp91_20 sp91_20 sp20_p3 11.551961
Rsn91_20 sn91_20 sn20_p3 11.551961
Rsp91_21 sp91_21 sp21_p3 11.551961
Rsn91_21 sn91_21 sn21_p3 11.551961
Rsp91_22 sp91_22 sp22_p3 11.551961
Rsn91_22 sn91_22 sn22_p3 11.551961
Rsp91_23 sp91_23 sp23_p3 11.551961
Rsn91_23 sn91_23 sn23_p3 11.551961
Rsp91_24 sp91_24 sp24_p3 11.551961
Rsn91_24 sn91_24 sn24_p3 11.551961
Rsp91_25 sp91_25 sp25_p3 11.551961
Rsn91_25 sn91_25 sn25_p3 11.551961
Rsp91_26 sp91_26 sp26_p3 11.551961
Rsn91_26 sn91_26 sn26_p3 11.551961
Rsp91_27 sp91_27 sp27_p3 11.551961
Rsn91_27 sn91_27 sn27_p3 11.551961
Rsp91_28 sp91_28 sp28_p3 11.551961
Rsn91_28 sn91_28 sn28_p3 11.551961
Rsp91_29 sp91_29 sp29_p3 11.551961
Rsn91_29 sn91_29 sn29_p3 11.551961
Rsp91_30 sp91_30 sp30_p3 11.551961
Rsn91_30 sn91_30 sn30_p3 11.551961
Rsp91_31 sp91_31 sp31_p3 11.551961
Rsn91_31 sn91_31 sn31_p3 11.551961
Rsp91_32 sp91_32 sp32_p3 11.551961
Rsn91_32 sn91_32 sn32_p3 11.551961
Rsp91_33 sp91_33 sp33_p3 11.551961
Rsn91_33 sn91_33 sn33_p3 11.551961
Rsp91_34 sp91_34 sp34_p3 11.551961
Rsn91_34 sn91_34 sn34_p3 11.551961
Rsp91_35 sp91_35 sp35_p3 11.551961
Rsn91_35 sn91_35 sn35_p3 11.551961
Rsp91_36 sp91_36 sp36_p3 11.551961
Rsn91_36 sn91_36 sn36_p3 11.551961
Rsp91_37 sp91_37 sp37_p3 11.551961
Rsn91_37 sn91_37 sn37_p3 11.551961
Rsp91_38 sp91_38 sp38_p3 11.551961
Rsn91_38 sn91_38 sn38_p3 11.551961
Rsp91_39 sp91_39 sp39_p3 11.551961
Rsn91_39 sn91_39 sn39_p3 11.551961
Rsp91_40 sp91_40 sp40_p3 11.551961
Rsn91_40 sn91_40 sn40_p3 11.551961
Rsp91_41 sp91_41 sp41_p3 11.551961
Rsn91_41 sn91_41 sn41_p3 11.551961
Rsp91_42 sp91_42 sp42_p3 11.551961
Rsn91_42 sn91_42 sn42_p3 11.551961
Rsp91_43 sp91_43 sp43_p3 11.551961
Rsn91_43 sn91_43 sn43_p3 11.551961
Rsp91_44 sp91_44 sp44_p3 11.551961
Rsn91_44 sn91_44 sn44_p3 11.551961
Rsp91_45 sp91_45 sp45_p3 11.551961
Rsn91_45 sn91_45 sn45_p3 11.551961
Rsp91_46 sp91_46 sp46_p3 11.551961
Rsn91_46 sn91_46 sn46_p3 11.551961
Rsp91_47 sp91_47 sp47_p3 11.551961
Rsn91_47 sn91_47 sn47_p3 11.551961
Rsp91_48 sp91_48 sp48_p3 11.551961
Rsn91_48 sn91_48 sn48_p3 11.551961
Rsp91_49 sp91_49 sp49_p3 11.551961
Rsn91_49 sn91_49 sn49_p3 11.551961
Rsp91_50 sp91_50 sp50_p3 11.551961
Rsn91_50 sn91_50 sn50_p3 11.551961
Rsp91_51 sp91_51 sp51_p3 11.551961
Rsn91_51 sn91_51 sn51_p3 11.551961
Rsp91_52 sp91_52 sp52_p3 11.551961
Rsn91_52 sn91_52 sn52_p3 11.551961
Rsp91_53 sp91_53 sp53_p3 11.551961
Rsn91_53 sn91_53 sn53_p3 11.551961
Rsp91_54 sp91_54 sp54_p3 11.551961
Rsn91_54 sn91_54 sn54_p3 11.551961
Rsp91_55 sp91_55 sp55_p3 11.551961
Rsn91_55 sn91_55 sn55_p3 11.551961
Rsp91_56 sp91_56 sp56_p3 11.551961
Rsn91_56 sn91_56 sn56_p3 11.551961
Rsp91_57 sp91_57 sp57_p3 11.551961
Rsn91_57 sn91_57 sn57_p3 11.551961
Rsp91_58 sp91_58 sp58_p3 11.551961
Rsn91_58 sn91_58 sn58_p3 11.551961
Rsp91_59 sp91_59 sp59_p3 11.551961
Rsn91_59 sn91_59 sn59_p3 11.551961
Rsp91_60 sp91_60 sp60_p3 11.551961
Rsn91_60 sn91_60 sn60_p3 11.551961
Rsp91_61 sp91_61 sp61_p3 11.551961
Rsn91_61 sn91_61 sn61_p3 11.551961
Rsp91_62 sp91_62 sp62_p3 11.551961
Rsn91_62 sn91_62 sn62_p3 11.551961
Rsp91_63 sp91_63 sp63_p3 11.551961
Rsn91_63 sn91_63 sn63_p3 11.551961
Rsp91_64 sp91_64 sp64_p3 11.551961
Rsn91_64 sn91_64 sn64_p3 11.551961
Rsp91_65 sp91_65 sp65_p3 11.551961
Rsn91_65 sn91_65 sn65_p3 11.551961
Rsp91_66 sp91_66 sp66_p3 11.551961
Rsn91_66 sn91_66 sn66_p3 11.551961
Rsp91_67 sp91_67 sp67_p3 11.551961
Rsn91_67 sn91_67 sn67_p3 11.551961
Rsp91_68 sp91_68 sp68_p3 11.551961
Rsn91_68 sn91_68 sn68_p3 11.551961
Rsp91_69 sp91_69 sp69_p3 11.551961
Rsn91_69 sn91_69 sn69_p3 11.551961
Rsp91_70 sp91_70 sp70_p3 11.551961
Rsn91_70 sn91_70 sn70_p3 11.551961
Rsp91_71 sp91_71 sp71_p3 11.551961
Rsn91_71 sn91_71 sn71_p3 11.551961
Rsp91_72 sp91_72 sp72_p3 11.551961
Rsn91_72 sn91_72 sn72_p3 11.551961
Rsp91_73 sp91_73 sp73_p3 11.551961
Rsn91_73 sn91_73 sn73_p3 11.551961
Rsp91_74 sp91_74 sp74_p3 11.551961
Rsn91_74 sn91_74 sn74_p3 11.551961
Rsp91_75 sp91_75 sp75_p3 11.551961
Rsn91_75 sn91_75 sn75_p3 11.551961
Rsp91_76 sp91_76 sp76_p3 11.551961
Rsn91_76 sn91_76 sn76_p3 11.551961
Rsp91_77 sp91_77 sp77_p3 11.551961
Rsn91_77 sn91_77 sn77_p3 11.551961
Rsp91_78 sp91_78 sp78_p3 11.551961
Rsn91_78 sn91_78 sn78_p3 11.551961
Rsp91_79 sp91_79 sp79_p3 11.551961
Rsn91_79 sn91_79 sn79_p3 11.551961
Rsp91_80 sp91_80 sp80_p3 11.551961
Rsn91_80 sn91_80 sn80_p3 11.551961
Rsp91_81 sp91_81 sp81_p3 11.551961
Rsn91_81 sn91_81 sn81_p3 11.551961
Rsp91_82 sp91_82 sp82_p3 11.551961
Rsn91_82 sn91_82 sn82_p3 11.551961
Rsp91_83 sp91_83 sp83_p3 11.551961
Rsn91_83 sn91_83 sn83_p3 11.551961
Rsp91_84 sp91_84 sp84_p3 11.551961
Rsn91_84 sn91_84 sn84_p3 11.551961
Rsp92_1 sp92_1 sp93_1 11.551961
Rsn92_1 sn92_1 sn93_1 11.551961
Rsp92_2 sp92_2 sp93_2 11.551961
Rsn92_2 sn92_2 sn93_2 11.551961
Rsp92_3 sp92_3 sp93_3 11.551961
Rsn92_3 sn92_3 sn93_3 11.551961
Rsp92_4 sp92_4 sp93_4 11.551961
Rsn92_4 sn92_4 sn93_4 11.551961
Rsp92_5 sp92_5 sp93_5 11.551961
Rsn92_5 sn92_5 sn93_5 11.551961
Rsp92_6 sp92_6 sp93_6 11.551961
Rsn92_6 sn92_6 sn93_6 11.551961
Rsp92_7 sp92_7 sp93_7 11.551961
Rsn92_7 sn92_7 sn93_7 11.551961
Rsp92_8 sp92_8 sp93_8 11.551961
Rsn92_8 sn92_8 sn93_8 11.551961
Rsp92_9 sp92_9 sp93_9 11.551961
Rsn92_9 sn92_9 sn93_9 11.551961
Rsp92_10 sp92_10 sp93_10 11.551961
Rsn92_10 sn92_10 sn93_10 11.551961
Rsp92_11 sp92_11 sp93_11 11.551961
Rsn92_11 sn92_11 sn93_11 11.551961
Rsp92_12 sp92_12 sp93_12 11.551961
Rsn92_12 sn92_12 sn93_12 11.551961
Rsp92_13 sp92_13 sp93_13 11.551961
Rsn92_13 sn92_13 sn93_13 11.551961
Rsp92_14 sp92_14 sp93_14 11.551961
Rsn92_14 sn92_14 sn93_14 11.551961
Rsp92_15 sp92_15 sp93_15 11.551961
Rsn92_15 sn92_15 sn93_15 11.551961
Rsp92_16 sp92_16 sp93_16 11.551961
Rsn92_16 sn92_16 sn93_16 11.551961
Rsp92_17 sp92_17 sp93_17 11.551961
Rsn92_17 sn92_17 sn93_17 11.551961
Rsp92_18 sp92_18 sp93_18 11.551961
Rsn92_18 sn92_18 sn93_18 11.551961
Rsp92_19 sp92_19 sp93_19 11.551961
Rsn92_19 sn92_19 sn93_19 11.551961
Rsp92_20 sp92_20 sp93_20 11.551961
Rsn92_20 sn92_20 sn93_20 11.551961
Rsp92_21 sp92_21 sp93_21 11.551961
Rsn92_21 sn92_21 sn93_21 11.551961
Rsp92_22 sp92_22 sp93_22 11.551961
Rsn92_22 sn92_22 sn93_22 11.551961
Rsp92_23 sp92_23 sp93_23 11.551961
Rsn92_23 sn92_23 sn93_23 11.551961
Rsp92_24 sp92_24 sp93_24 11.551961
Rsn92_24 sn92_24 sn93_24 11.551961
Rsp92_25 sp92_25 sp93_25 11.551961
Rsn92_25 sn92_25 sn93_25 11.551961
Rsp92_26 sp92_26 sp93_26 11.551961
Rsn92_26 sn92_26 sn93_26 11.551961
Rsp92_27 sp92_27 sp93_27 11.551961
Rsn92_27 sn92_27 sn93_27 11.551961
Rsp92_28 sp92_28 sp93_28 11.551961
Rsn92_28 sn92_28 sn93_28 11.551961
Rsp92_29 sp92_29 sp93_29 11.551961
Rsn92_29 sn92_29 sn93_29 11.551961
Rsp92_30 sp92_30 sp93_30 11.551961
Rsn92_30 sn92_30 sn93_30 11.551961
Rsp92_31 sp92_31 sp93_31 11.551961
Rsn92_31 sn92_31 sn93_31 11.551961
Rsp92_32 sp92_32 sp93_32 11.551961
Rsn92_32 sn92_32 sn93_32 11.551961
Rsp92_33 sp92_33 sp93_33 11.551961
Rsn92_33 sn92_33 sn93_33 11.551961
Rsp92_34 sp92_34 sp93_34 11.551961
Rsn92_34 sn92_34 sn93_34 11.551961
Rsp92_35 sp92_35 sp93_35 11.551961
Rsn92_35 sn92_35 sn93_35 11.551961
Rsp92_36 sp92_36 sp93_36 11.551961
Rsn92_36 sn92_36 sn93_36 11.551961
Rsp92_37 sp92_37 sp93_37 11.551961
Rsn92_37 sn92_37 sn93_37 11.551961
Rsp92_38 sp92_38 sp93_38 11.551961
Rsn92_38 sn92_38 sn93_38 11.551961
Rsp92_39 sp92_39 sp93_39 11.551961
Rsn92_39 sn92_39 sn93_39 11.551961
Rsp92_40 sp92_40 sp93_40 11.551961
Rsn92_40 sn92_40 sn93_40 11.551961
Rsp92_41 sp92_41 sp93_41 11.551961
Rsn92_41 sn92_41 sn93_41 11.551961
Rsp92_42 sp92_42 sp93_42 11.551961
Rsn92_42 sn92_42 sn93_42 11.551961
Rsp92_43 sp92_43 sp93_43 11.551961
Rsn92_43 sn92_43 sn93_43 11.551961
Rsp92_44 sp92_44 sp93_44 11.551961
Rsn92_44 sn92_44 sn93_44 11.551961
Rsp92_45 sp92_45 sp93_45 11.551961
Rsn92_45 sn92_45 sn93_45 11.551961
Rsp92_46 sp92_46 sp93_46 11.551961
Rsn92_46 sn92_46 sn93_46 11.551961
Rsp92_47 sp92_47 sp93_47 11.551961
Rsn92_47 sn92_47 sn93_47 11.551961
Rsp92_48 sp92_48 sp93_48 11.551961
Rsn92_48 sn92_48 sn93_48 11.551961
Rsp92_49 sp92_49 sp93_49 11.551961
Rsn92_49 sn92_49 sn93_49 11.551961
Rsp92_50 sp92_50 sp93_50 11.551961
Rsn92_50 sn92_50 sn93_50 11.551961
Rsp92_51 sp92_51 sp93_51 11.551961
Rsn92_51 sn92_51 sn93_51 11.551961
Rsp92_52 sp92_52 sp93_52 11.551961
Rsn92_52 sn92_52 sn93_52 11.551961
Rsp92_53 sp92_53 sp93_53 11.551961
Rsn92_53 sn92_53 sn93_53 11.551961
Rsp92_54 sp92_54 sp93_54 11.551961
Rsn92_54 sn92_54 sn93_54 11.551961
Rsp92_55 sp92_55 sp93_55 11.551961
Rsn92_55 sn92_55 sn93_55 11.551961
Rsp92_56 sp92_56 sp93_56 11.551961
Rsn92_56 sn92_56 sn93_56 11.551961
Rsp92_57 sp92_57 sp93_57 11.551961
Rsn92_57 sn92_57 sn93_57 11.551961
Rsp92_58 sp92_58 sp93_58 11.551961
Rsn92_58 sn92_58 sn93_58 11.551961
Rsp92_59 sp92_59 sp93_59 11.551961
Rsn92_59 sn92_59 sn93_59 11.551961
Rsp92_60 sp92_60 sp93_60 11.551961
Rsn92_60 sn92_60 sn93_60 11.551961
Rsp92_61 sp92_61 sp93_61 11.551961
Rsn92_61 sn92_61 sn93_61 11.551961
Rsp92_62 sp92_62 sp93_62 11.551961
Rsn92_62 sn92_62 sn93_62 11.551961
Rsp92_63 sp92_63 sp93_63 11.551961
Rsn92_63 sn92_63 sn93_63 11.551961
Rsp92_64 sp92_64 sp93_64 11.551961
Rsn92_64 sn92_64 sn93_64 11.551961
Rsp92_65 sp92_65 sp93_65 11.551961
Rsn92_65 sn92_65 sn93_65 11.551961
Rsp92_66 sp92_66 sp93_66 11.551961
Rsn92_66 sn92_66 sn93_66 11.551961
Rsp92_67 sp92_67 sp93_67 11.551961
Rsn92_67 sn92_67 sn93_67 11.551961
Rsp92_68 sp92_68 sp93_68 11.551961
Rsn92_68 sn92_68 sn93_68 11.551961
Rsp92_69 sp92_69 sp93_69 11.551961
Rsn92_69 sn92_69 sn93_69 11.551961
Rsp92_70 sp92_70 sp93_70 11.551961
Rsn92_70 sn92_70 sn93_70 11.551961
Rsp92_71 sp92_71 sp93_71 11.551961
Rsn92_71 sn92_71 sn93_71 11.551961
Rsp92_72 sp92_72 sp93_72 11.551961
Rsn92_72 sn92_72 sn93_72 11.551961
Rsp92_73 sp92_73 sp93_73 11.551961
Rsn92_73 sn92_73 sn93_73 11.551961
Rsp92_74 sp92_74 sp93_74 11.551961
Rsn92_74 sn92_74 sn93_74 11.551961
Rsp92_75 sp92_75 sp93_75 11.551961
Rsn92_75 sn92_75 sn93_75 11.551961
Rsp92_76 sp92_76 sp93_76 11.551961
Rsn92_76 sn92_76 sn93_76 11.551961
Rsp92_77 sp92_77 sp93_77 11.551961
Rsn92_77 sn92_77 sn93_77 11.551961
Rsp92_78 sp92_78 sp93_78 11.551961
Rsn92_78 sn92_78 sn93_78 11.551961
Rsp92_79 sp92_79 sp93_79 11.551961
Rsn92_79 sn92_79 sn93_79 11.551961
Rsp92_80 sp92_80 sp93_80 11.551961
Rsn92_80 sn92_80 sn93_80 11.551961
Rsp92_81 sp92_81 sp93_81 11.551961
Rsn92_81 sn92_81 sn93_81 11.551961
Rsp92_82 sp92_82 sp93_82 11.551961
Rsn92_82 sn92_82 sn93_82 11.551961
Rsp92_83 sp92_83 sp93_83 11.551961
Rsn92_83 sn92_83 sn93_83 11.551961
Rsp92_84 sp92_84 sp93_84 11.551961
Rsn92_84 sn92_84 sn93_84 11.551961
Rsp93_1 sp93_1 sp94_1 11.551961
Rsn93_1 sn93_1 sn94_1 11.551961
Rsp93_2 sp93_2 sp94_2 11.551961
Rsn93_2 sn93_2 sn94_2 11.551961
Rsp93_3 sp93_3 sp94_3 11.551961
Rsn93_3 sn93_3 sn94_3 11.551961
Rsp93_4 sp93_4 sp94_4 11.551961
Rsn93_4 sn93_4 sn94_4 11.551961
Rsp93_5 sp93_5 sp94_5 11.551961
Rsn93_5 sn93_5 sn94_5 11.551961
Rsp93_6 sp93_6 sp94_6 11.551961
Rsn93_6 sn93_6 sn94_6 11.551961
Rsp93_7 sp93_7 sp94_7 11.551961
Rsn93_7 sn93_7 sn94_7 11.551961
Rsp93_8 sp93_8 sp94_8 11.551961
Rsn93_8 sn93_8 sn94_8 11.551961
Rsp93_9 sp93_9 sp94_9 11.551961
Rsn93_9 sn93_9 sn94_9 11.551961
Rsp93_10 sp93_10 sp94_10 11.551961
Rsn93_10 sn93_10 sn94_10 11.551961
Rsp93_11 sp93_11 sp94_11 11.551961
Rsn93_11 sn93_11 sn94_11 11.551961
Rsp93_12 sp93_12 sp94_12 11.551961
Rsn93_12 sn93_12 sn94_12 11.551961
Rsp93_13 sp93_13 sp94_13 11.551961
Rsn93_13 sn93_13 sn94_13 11.551961
Rsp93_14 sp93_14 sp94_14 11.551961
Rsn93_14 sn93_14 sn94_14 11.551961
Rsp93_15 sp93_15 sp94_15 11.551961
Rsn93_15 sn93_15 sn94_15 11.551961
Rsp93_16 sp93_16 sp94_16 11.551961
Rsn93_16 sn93_16 sn94_16 11.551961
Rsp93_17 sp93_17 sp94_17 11.551961
Rsn93_17 sn93_17 sn94_17 11.551961
Rsp93_18 sp93_18 sp94_18 11.551961
Rsn93_18 sn93_18 sn94_18 11.551961
Rsp93_19 sp93_19 sp94_19 11.551961
Rsn93_19 sn93_19 sn94_19 11.551961
Rsp93_20 sp93_20 sp94_20 11.551961
Rsn93_20 sn93_20 sn94_20 11.551961
Rsp93_21 sp93_21 sp94_21 11.551961
Rsn93_21 sn93_21 sn94_21 11.551961
Rsp93_22 sp93_22 sp94_22 11.551961
Rsn93_22 sn93_22 sn94_22 11.551961
Rsp93_23 sp93_23 sp94_23 11.551961
Rsn93_23 sn93_23 sn94_23 11.551961
Rsp93_24 sp93_24 sp94_24 11.551961
Rsn93_24 sn93_24 sn94_24 11.551961
Rsp93_25 sp93_25 sp94_25 11.551961
Rsn93_25 sn93_25 sn94_25 11.551961
Rsp93_26 sp93_26 sp94_26 11.551961
Rsn93_26 sn93_26 sn94_26 11.551961
Rsp93_27 sp93_27 sp94_27 11.551961
Rsn93_27 sn93_27 sn94_27 11.551961
Rsp93_28 sp93_28 sp94_28 11.551961
Rsn93_28 sn93_28 sn94_28 11.551961
Rsp93_29 sp93_29 sp94_29 11.551961
Rsn93_29 sn93_29 sn94_29 11.551961
Rsp93_30 sp93_30 sp94_30 11.551961
Rsn93_30 sn93_30 sn94_30 11.551961
Rsp93_31 sp93_31 sp94_31 11.551961
Rsn93_31 sn93_31 sn94_31 11.551961
Rsp93_32 sp93_32 sp94_32 11.551961
Rsn93_32 sn93_32 sn94_32 11.551961
Rsp93_33 sp93_33 sp94_33 11.551961
Rsn93_33 sn93_33 sn94_33 11.551961
Rsp93_34 sp93_34 sp94_34 11.551961
Rsn93_34 sn93_34 sn94_34 11.551961
Rsp93_35 sp93_35 sp94_35 11.551961
Rsn93_35 sn93_35 sn94_35 11.551961
Rsp93_36 sp93_36 sp94_36 11.551961
Rsn93_36 sn93_36 sn94_36 11.551961
Rsp93_37 sp93_37 sp94_37 11.551961
Rsn93_37 sn93_37 sn94_37 11.551961
Rsp93_38 sp93_38 sp94_38 11.551961
Rsn93_38 sn93_38 sn94_38 11.551961
Rsp93_39 sp93_39 sp94_39 11.551961
Rsn93_39 sn93_39 sn94_39 11.551961
Rsp93_40 sp93_40 sp94_40 11.551961
Rsn93_40 sn93_40 sn94_40 11.551961
Rsp93_41 sp93_41 sp94_41 11.551961
Rsn93_41 sn93_41 sn94_41 11.551961
Rsp93_42 sp93_42 sp94_42 11.551961
Rsn93_42 sn93_42 sn94_42 11.551961
Rsp93_43 sp93_43 sp94_43 11.551961
Rsn93_43 sn93_43 sn94_43 11.551961
Rsp93_44 sp93_44 sp94_44 11.551961
Rsn93_44 sn93_44 sn94_44 11.551961
Rsp93_45 sp93_45 sp94_45 11.551961
Rsn93_45 sn93_45 sn94_45 11.551961
Rsp93_46 sp93_46 sp94_46 11.551961
Rsn93_46 sn93_46 sn94_46 11.551961
Rsp93_47 sp93_47 sp94_47 11.551961
Rsn93_47 sn93_47 sn94_47 11.551961
Rsp93_48 sp93_48 sp94_48 11.551961
Rsn93_48 sn93_48 sn94_48 11.551961
Rsp93_49 sp93_49 sp94_49 11.551961
Rsn93_49 sn93_49 sn94_49 11.551961
Rsp93_50 sp93_50 sp94_50 11.551961
Rsn93_50 sn93_50 sn94_50 11.551961
Rsp93_51 sp93_51 sp94_51 11.551961
Rsn93_51 sn93_51 sn94_51 11.551961
Rsp93_52 sp93_52 sp94_52 11.551961
Rsn93_52 sn93_52 sn94_52 11.551961
Rsp93_53 sp93_53 sp94_53 11.551961
Rsn93_53 sn93_53 sn94_53 11.551961
Rsp93_54 sp93_54 sp94_54 11.551961
Rsn93_54 sn93_54 sn94_54 11.551961
Rsp93_55 sp93_55 sp94_55 11.551961
Rsn93_55 sn93_55 sn94_55 11.551961
Rsp93_56 sp93_56 sp94_56 11.551961
Rsn93_56 sn93_56 sn94_56 11.551961
Rsp93_57 sp93_57 sp94_57 11.551961
Rsn93_57 sn93_57 sn94_57 11.551961
Rsp93_58 sp93_58 sp94_58 11.551961
Rsn93_58 sn93_58 sn94_58 11.551961
Rsp93_59 sp93_59 sp94_59 11.551961
Rsn93_59 sn93_59 sn94_59 11.551961
Rsp93_60 sp93_60 sp94_60 11.551961
Rsn93_60 sn93_60 sn94_60 11.551961
Rsp93_61 sp93_61 sp94_61 11.551961
Rsn93_61 sn93_61 sn94_61 11.551961
Rsp93_62 sp93_62 sp94_62 11.551961
Rsn93_62 sn93_62 sn94_62 11.551961
Rsp93_63 sp93_63 sp94_63 11.551961
Rsn93_63 sn93_63 sn94_63 11.551961
Rsp93_64 sp93_64 sp94_64 11.551961
Rsn93_64 sn93_64 sn94_64 11.551961
Rsp93_65 sp93_65 sp94_65 11.551961
Rsn93_65 sn93_65 sn94_65 11.551961
Rsp93_66 sp93_66 sp94_66 11.551961
Rsn93_66 sn93_66 sn94_66 11.551961
Rsp93_67 sp93_67 sp94_67 11.551961
Rsn93_67 sn93_67 sn94_67 11.551961
Rsp93_68 sp93_68 sp94_68 11.551961
Rsn93_68 sn93_68 sn94_68 11.551961
Rsp93_69 sp93_69 sp94_69 11.551961
Rsn93_69 sn93_69 sn94_69 11.551961
Rsp93_70 sp93_70 sp94_70 11.551961
Rsn93_70 sn93_70 sn94_70 11.551961
Rsp93_71 sp93_71 sp94_71 11.551961
Rsn93_71 sn93_71 sn94_71 11.551961
Rsp93_72 sp93_72 sp94_72 11.551961
Rsn93_72 sn93_72 sn94_72 11.551961
Rsp93_73 sp93_73 sp94_73 11.551961
Rsn93_73 sn93_73 sn94_73 11.551961
Rsp93_74 sp93_74 sp94_74 11.551961
Rsn93_74 sn93_74 sn94_74 11.551961
Rsp93_75 sp93_75 sp94_75 11.551961
Rsn93_75 sn93_75 sn94_75 11.551961
Rsp93_76 sp93_76 sp94_76 11.551961
Rsn93_76 sn93_76 sn94_76 11.551961
Rsp93_77 sp93_77 sp94_77 11.551961
Rsn93_77 sn93_77 sn94_77 11.551961
Rsp93_78 sp93_78 sp94_78 11.551961
Rsn93_78 sn93_78 sn94_78 11.551961
Rsp93_79 sp93_79 sp94_79 11.551961
Rsn93_79 sn93_79 sn94_79 11.551961
Rsp93_80 sp93_80 sp94_80 11.551961
Rsn93_80 sn93_80 sn94_80 11.551961
Rsp93_81 sp93_81 sp94_81 11.551961
Rsn93_81 sn93_81 sn94_81 11.551961
Rsp93_82 sp93_82 sp94_82 11.551961
Rsn93_82 sn93_82 sn94_82 11.551961
Rsp93_83 sp93_83 sp94_83 11.551961
Rsn93_83 sn93_83 sn94_83 11.551961
Rsp93_84 sp93_84 sp94_84 11.551961
Rsn93_84 sn93_84 sn94_84 11.551961
Rsp94_1 sp94_1 sp95_1 11.551961
Rsn94_1 sn94_1 sn95_1 11.551961
Rsp94_2 sp94_2 sp95_2 11.551961
Rsn94_2 sn94_2 sn95_2 11.551961
Rsp94_3 sp94_3 sp95_3 11.551961
Rsn94_3 sn94_3 sn95_3 11.551961
Rsp94_4 sp94_4 sp95_4 11.551961
Rsn94_4 sn94_4 sn95_4 11.551961
Rsp94_5 sp94_5 sp95_5 11.551961
Rsn94_5 sn94_5 sn95_5 11.551961
Rsp94_6 sp94_6 sp95_6 11.551961
Rsn94_6 sn94_6 sn95_6 11.551961
Rsp94_7 sp94_7 sp95_7 11.551961
Rsn94_7 sn94_7 sn95_7 11.551961
Rsp94_8 sp94_8 sp95_8 11.551961
Rsn94_8 sn94_8 sn95_8 11.551961
Rsp94_9 sp94_9 sp95_9 11.551961
Rsn94_9 sn94_9 sn95_9 11.551961
Rsp94_10 sp94_10 sp95_10 11.551961
Rsn94_10 sn94_10 sn95_10 11.551961
Rsp94_11 sp94_11 sp95_11 11.551961
Rsn94_11 sn94_11 sn95_11 11.551961
Rsp94_12 sp94_12 sp95_12 11.551961
Rsn94_12 sn94_12 sn95_12 11.551961
Rsp94_13 sp94_13 sp95_13 11.551961
Rsn94_13 sn94_13 sn95_13 11.551961
Rsp94_14 sp94_14 sp95_14 11.551961
Rsn94_14 sn94_14 sn95_14 11.551961
Rsp94_15 sp94_15 sp95_15 11.551961
Rsn94_15 sn94_15 sn95_15 11.551961
Rsp94_16 sp94_16 sp95_16 11.551961
Rsn94_16 sn94_16 sn95_16 11.551961
Rsp94_17 sp94_17 sp95_17 11.551961
Rsn94_17 sn94_17 sn95_17 11.551961
Rsp94_18 sp94_18 sp95_18 11.551961
Rsn94_18 sn94_18 sn95_18 11.551961
Rsp94_19 sp94_19 sp95_19 11.551961
Rsn94_19 sn94_19 sn95_19 11.551961
Rsp94_20 sp94_20 sp95_20 11.551961
Rsn94_20 sn94_20 sn95_20 11.551961
Rsp94_21 sp94_21 sp95_21 11.551961
Rsn94_21 sn94_21 sn95_21 11.551961
Rsp94_22 sp94_22 sp95_22 11.551961
Rsn94_22 sn94_22 sn95_22 11.551961
Rsp94_23 sp94_23 sp95_23 11.551961
Rsn94_23 sn94_23 sn95_23 11.551961
Rsp94_24 sp94_24 sp95_24 11.551961
Rsn94_24 sn94_24 sn95_24 11.551961
Rsp94_25 sp94_25 sp95_25 11.551961
Rsn94_25 sn94_25 sn95_25 11.551961
Rsp94_26 sp94_26 sp95_26 11.551961
Rsn94_26 sn94_26 sn95_26 11.551961
Rsp94_27 sp94_27 sp95_27 11.551961
Rsn94_27 sn94_27 sn95_27 11.551961
Rsp94_28 sp94_28 sp95_28 11.551961
Rsn94_28 sn94_28 sn95_28 11.551961
Rsp94_29 sp94_29 sp95_29 11.551961
Rsn94_29 sn94_29 sn95_29 11.551961
Rsp94_30 sp94_30 sp95_30 11.551961
Rsn94_30 sn94_30 sn95_30 11.551961
Rsp94_31 sp94_31 sp95_31 11.551961
Rsn94_31 sn94_31 sn95_31 11.551961
Rsp94_32 sp94_32 sp95_32 11.551961
Rsn94_32 sn94_32 sn95_32 11.551961
Rsp94_33 sp94_33 sp95_33 11.551961
Rsn94_33 sn94_33 sn95_33 11.551961
Rsp94_34 sp94_34 sp95_34 11.551961
Rsn94_34 sn94_34 sn95_34 11.551961
Rsp94_35 sp94_35 sp95_35 11.551961
Rsn94_35 sn94_35 sn95_35 11.551961
Rsp94_36 sp94_36 sp95_36 11.551961
Rsn94_36 sn94_36 sn95_36 11.551961
Rsp94_37 sp94_37 sp95_37 11.551961
Rsn94_37 sn94_37 sn95_37 11.551961
Rsp94_38 sp94_38 sp95_38 11.551961
Rsn94_38 sn94_38 sn95_38 11.551961
Rsp94_39 sp94_39 sp95_39 11.551961
Rsn94_39 sn94_39 sn95_39 11.551961
Rsp94_40 sp94_40 sp95_40 11.551961
Rsn94_40 sn94_40 sn95_40 11.551961
Rsp94_41 sp94_41 sp95_41 11.551961
Rsn94_41 sn94_41 sn95_41 11.551961
Rsp94_42 sp94_42 sp95_42 11.551961
Rsn94_42 sn94_42 sn95_42 11.551961
Rsp94_43 sp94_43 sp95_43 11.551961
Rsn94_43 sn94_43 sn95_43 11.551961
Rsp94_44 sp94_44 sp95_44 11.551961
Rsn94_44 sn94_44 sn95_44 11.551961
Rsp94_45 sp94_45 sp95_45 11.551961
Rsn94_45 sn94_45 sn95_45 11.551961
Rsp94_46 sp94_46 sp95_46 11.551961
Rsn94_46 sn94_46 sn95_46 11.551961
Rsp94_47 sp94_47 sp95_47 11.551961
Rsn94_47 sn94_47 sn95_47 11.551961
Rsp94_48 sp94_48 sp95_48 11.551961
Rsn94_48 sn94_48 sn95_48 11.551961
Rsp94_49 sp94_49 sp95_49 11.551961
Rsn94_49 sn94_49 sn95_49 11.551961
Rsp94_50 sp94_50 sp95_50 11.551961
Rsn94_50 sn94_50 sn95_50 11.551961
Rsp94_51 sp94_51 sp95_51 11.551961
Rsn94_51 sn94_51 sn95_51 11.551961
Rsp94_52 sp94_52 sp95_52 11.551961
Rsn94_52 sn94_52 sn95_52 11.551961
Rsp94_53 sp94_53 sp95_53 11.551961
Rsn94_53 sn94_53 sn95_53 11.551961
Rsp94_54 sp94_54 sp95_54 11.551961
Rsn94_54 sn94_54 sn95_54 11.551961
Rsp94_55 sp94_55 sp95_55 11.551961
Rsn94_55 sn94_55 sn95_55 11.551961
Rsp94_56 sp94_56 sp95_56 11.551961
Rsn94_56 sn94_56 sn95_56 11.551961
Rsp94_57 sp94_57 sp95_57 11.551961
Rsn94_57 sn94_57 sn95_57 11.551961
Rsp94_58 sp94_58 sp95_58 11.551961
Rsn94_58 sn94_58 sn95_58 11.551961
Rsp94_59 sp94_59 sp95_59 11.551961
Rsn94_59 sn94_59 sn95_59 11.551961
Rsp94_60 sp94_60 sp95_60 11.551961
Rsn94_60 sn94_60 sn95_60 11.551961
Rsp94_61 sp94_61 sp95_61 11.551961
Rsn94_61 sn94_61 sn95_61 11.551961
Rsp94_62 sp94_62 sp95_62 11.551961
Rsn94_62 sn94_62 sn95_62 11.551961
Rsp94_63 sp94_63 sp95_63 11.551961
Rsn94_63 sn94_63 sn95_63 11.551961
Rsp94_64 sp94_64 sp95_64 11.551961
Rsn94_64 sn94_64 sn95_64 11.551961
Rsp94_65 sp94_65 sp95_65 11.551961
Rsn94_65 sn94_65 sn95_65 11.551961
Rsp94_66 sp94_66 sp95_66 11.551961
Rsn94_66 sn94_66 sn95_66 11.551961
Rsp94_67 sp94_67 sp95_67 11.551961
Rsn94_67 sn94_67 sn95_67 11.551961
Rsp94_68 sp94_68 sp95_68 11.551961
Rsn94_68 sn94_68 sn95_68 11.551961
Rsp94_69 sp94_69 sp95_69 11.551961
Rsn94_69 sn94_69 sn95_69 11.551961
Rsp94_70 sp94_70 sp95_70 11.551961
Rsn94_70 sn94_70 sn95_70 11.551961
Rsp94_71 sp94_71 sp95_71 11.551961
Rsn94_71 sn94_71 sn95_71 11.551961
Rsp94_72 sp94_72 sp95_72 11.551961
Rsn94_72 sn94_72 sn95_72 11.551961
Rsp94_73 sp94_73 sp95_73 11.551961
Rsn94_73 sn94_73 sn95_73 11.551961
Rsp94_74 sp94_74 sp95_74 11.551961
Rsn94_74 sn94_74 sn95_74 11.551961
Rsp94_75 sp94_75 sp95_75 11.551961
Rsn94_75 sn94_75 sn95_75 11.551961
Rsp94_76 sp94_76 sp95_76 11.551961
Rsn94_76 sn94_76 sn95_76 11.551961
Rsp94_77 sp94_77 sp95_77 11.551961
Rsn94_77 sn94_77 sn95_77 11.551961
Rsp94_78 sp94_78 sp95_78 11.551961
Rsn94_78 sn94_78 sn95_78 11.551961
Rsp94_79 sp94_79 sp95_79 11.551961
Rsn94_79 sn94_79 sn95_79 11.551961
Rsp94_80 sp94_80 sp95_80 11.551961
Rsn94_80 sn94_80 sn95_80 11.551961
Rsp94_81 sp94_81 sp95_81 11.551961
Rsn94_81 sn94_81 sn95_81 11.551961
Rsp94_82 sp94_82 sp95_82 11.551961
Rsn94_82 sn94_82 sn95_82 11.551961
Rsp94_83 sp94_83 sp95_83 11.551961
Rsn94_83 sn94_83 sn95_83 11.551961
Rsp94_84 sp94_84 sp95_84 11.551961
Rsn94_84 sn94_84 sn95_84 11.551961
Rsp95_1 sp95_1 sp96_1 11.551961
Rsn95_1 sn95_1 sn96_1 11.551961
Rsp95_2 sp95_2 sp96_2 11.551961
Rsn95_2 sn95_2 sn96_2 11.551961
Rsp95_3 sp95_3 sp96_3 11.551961
Rsn95_3 sn95_3 sn96_3 11.551961
Rsp95_4 sp95_4 sp96_4 11.551961
Rsn95_4 sn95_4 sn96_4 11.551961
Rsp95_5 sp95_5 sp96_5 11.551961
Rsn95_5 sn95_5 sn96_5 11.551961
Rsp95_6 sp95_6 sp96_6 11.551961
Rsn95_6 sn95_6 sn96_6 11.551961
Rsp95_7 sp95_7 sp96_7 11.551961
Rsn95_7 sn95_7 sn96_7 11.551961
Rsp95_8 sp95_8 sp96_8 11.551961
Rsn95_8 sn95_8 sn96_8 11.551961
Rsp95_9 sp95_9 sp96_9 11.551961
Rsn95_9 sn95_9 sn96_9 11.551961
Rsp95_10 sp95_10 sp96_10 11.551961
Rsn95_10 sn95_10 sn96_10 11.551961
Rsp95_11 sp95_11 sp96_11 11.551961
Rsn95_11 sn95_11 sn96_11 11.551961
Rsp95_12 sp95_12 sp96_12 11.551961
Rsn95_12 sn95_12 sn96_12 11.551961
Rsp95_13 sp95_13 sp96_13 11.551961
Rsn95_13 sn95_13 sn96_13 11.551961
Rsp95_14 sp95_14 sp96_14 11.551961
Rsn95_14 sn95_14 sn96_14 11.551961
Rsp95_15 sp95_15 sp96_15 11.551961
Rsn95_15 sn95_15 sn96_15 11.551961
Rsp95_16 sp95_16 sp96_16 11.551961
Rsn95_16 sn95_16 sn96_16 11.551961
Rsp95_17 sp95_17 sp96_17 11.551961
Rsn95_17 sn95_17 sn96_17 11.551961
Rsp95_18 sp95_18 sp96_18 11.551961
Rsn95_18 sn95_18 sn96_18 11.551961
Rsp95_19 sp95_19 sp96_19 11.551961
Rsn95_19 sn95_19 sn96_19 11.551961
Rsp95_20 sp95_20 sp96_20 11.551961
Rsn95_20 sn95_20 sn96_20 11.551961
Rsp95_21 sp95_21 sp96_21 11.551961
Rsn95_21 sn95_21 sn96_21 11.551961
Rsp95_22 sp95_22 sp96_22 11.551961
Rsn95_22 sn95_22 sn96_22 11.551961
Rsp95_23 sp95_23 sp96_23 11.551961
Rsn95_23 sn95_23 sn96_23 11.551961
Rsp95_24 sp95_24 sp96_24 11.551961
Rsn95_24 sn95_24 sn96_24 11.551961
Rsp95_25 sp95_25 sp96_25 11.551961
Rsn95_25 sn95_25 sn96_25 11.551961
Rsp95_26 sp95_26 sp96_26 11.551961
Rsn95_26 sn95_26 sn96_26 11.551961
Rsp95_27 sp95_27 sp96_27 11.551961
Rsn95_27 sn95_27 sn96_27 11.551961
Rsp95_28 sp95_28 sp96_28 11.551961
Rsn95_28 sn95_28 sn96_28 11.551961
Rsp95_29 sp95_29 sp96_29 11.551961
Rsn95_29 sn95_29 sn96_29 11.551961
Rsp95_30 sp95_30 sp96_30 11.551961
Rsn95_30 sn95_30 sn96_30 11.551961
Rsp95_31 sp95_31 sp96_31 11.551961
Rsn95_31 sn95_31 sn96_31 11.551961
Rsp95_32 sp95_32 sp96_32 11.551961
Rsn95_32 sn95_32 sn96_32 11.551961
Rsp95_33 sp95_33 sp96_33 11.551961
Rsn95_33 sn95_33 sn96_33 11.551961
Rsp95_34 sp95_34 sp96_34 11.551961
Rsn95_34 sn95_34 sn96_34 11.551961
Rsp95_35 sp95_35 sp96_35 11.551961
Rsn95_35 sn95_35 sn96_35 11.551961
Rsp95_36 sp95_36 sp96_36 11.551961
Rsn95_36 sn95_36 sn96_36 11.551961
Rsp95_37 sp95_37 sp96_37 11.551961
Rsn95_37 sn95_37 sn96_37 11.551961
Rsp95_38 sp95_38 sp96_38 11.551961
Rsn95_38 sn95_38 sn96_38 11.551961
Rsp95_39 sp95_39 sp96_39 11.551961
Rsn95_39 sn95_39 sn96_39 11.551961
Rsp95_40 sp95_40 sp96_40 11.551961
Rsn95_40 sn95_40 sn96_40 11.551961
Rsp95_41 sp95_41 sp96_41 11.551961
Rsn95_41 sn95_41 sn96_41 11.551961
Rsp95_42 sp95_42 sp96_42 11.551961
Rsn95_42 sn95_42 sn96_42 11.551961
Rsp95_43 sp95_43 sp96_43 11.551961
Rsn95_43 sn95_43 sn96_43 11.551961
Rsp95_44 sp95_44 sp96_44 11.551961
Rsn95_44 sn95_44 sn96_44 11.551961
Rsp95_45 sp95_45 sp96_45 11.551961
Rsn95_45 sn95_45 sn96_45 11.551961
Rsp95_46 sp95_46 sp96_46 11.551961
Rsn95_46 sn95_46 sn96_46 11.551961
Rsp95_47 sp95_47 sp96_47 11.551961
Rsn95_47 sn95_47 sn96_47 11.551961
Rsp95_48 sp95_48 sp96_48 11.551961
Rsn95_48 sn95_48 sn96_48 11.551961
Rsp95_49 sp95_49 sp96_49 11.551961
Rsn95_49 sn95_49 sn96_49 11.551961
Rsp95_50 sp95_50 sp96_50 11.551961
Rsn95_50 sn95_50 sn96_50 11.551961
Rsp95_51 sp95_51 sp96_51 11.551961
Rsn95_51 sn95_51 sn96_51 11.551961
Rsp95_52 sp95_52 sp96_52 11.551961
Rsn95_52 sn95_52 sn96_52 11.551961
Rsp95_53 sp95_53 sp96_53 11.551961
Rsn95_53 sn95_53 sn96_53 11.551961
Rsp95_54 sp95_54 sp96_54 11.551961
Rsn95_54 sn95_54 sn96_54 11.551961
Rsp95_55 sp95_55 sp96_55 11.551961
Rsn95_55 sn95_55 sn96_55 11.551961
Rsp95_56 sp95_56 sp96_56 11.551961
Rsn95_56 sn95_56 sn96_56 11.551961
Rsp95_57 sp95_57 sp96_57 11.551961
Rsn95_57 sn95_57 sn96_57 11.551961
Rsp95_58 sp95_58 sp96_58 11.551961
Rsn95_58 sn95_58 sn96_58 11.551961
Rsp95_59 sp95_59 sp96_59 11.551961
Rsn95_59 sn95_59 sn96_59 11.551961
Rsp95_60 sp95_60 sp96_60 11.551961
Rsn95_60 sn95_60 sn96_60 11.551961
Rsp95_61 sp95_61 sp96_61 11.551961
Rsn95_61 sn95_61 sn96_61 11.551961
Rsp95_62 sp95_62 sp96_62 11.551961
Rsn95_62 sn95_62 sn96_62 11.551961
Rsp95_63 sp95_63 sp96_63 11.551961
Rsn95_63 sn95_63 sn96_63 11.551961
Rsp95_64 sp95_64 sp96_64 11.551961
Rsn95_64 sn95_64 sn96_64 11.551961
Rsp95_65 sp95_65 sp96_65 11.551961
Rsn95_65 sn95_65 sn96_65 11.551961
Rsp95_66 sp95_66 sp96_66 11.551961
Rsn95_66 sn95_66 sn96_66 11.551961
Rsp95_67 sp95_67 sp96_67 11.551961
Rsn95_67 sn95_67 sn96_67 11.551961
Rsp95_68 sp95_68 sp96_68 11.551961
Rsn95_68 sn95_68 sn96_68 11.551961
Rsp95_69 sp95_69 sp96_69 11.551961
Rsn95_69 sn95_69 sn96_69 11.551961
Rsp95_70 sp95_70 sp96_70 11.551961
Rsn95_70 sn95_70 sn96_70 11.551961
Rsp95_71 sp95_71 sp96_71 11.551961
Rsn95_71 sn95_71 sn96_71 11.551961
Rsp95_72 sp95_72 sp96_72 11.551961
Rsn95_72 sn95_72 sn96_72 11.551961
Rsp95_73 sp95_73 sp96_73 11.551961
Rsn95_73 sn95_73 sn96_73 11.551961
Rsp95_74 sp95_74 sp96_74 11.551961
Rsn95_74 sn95_74 sn96_74 11.551961
Rsp95_75 sp95_75 sp96_75 11.551961
Rsn95_75 sn95_75 sn96_75 11.551961
Rsp95_76 sp95_76 sp96_76 11.551961
Rsn95_76 sn95_76 sn96_76 11.551961
Rsp95_77 sp95_77 sp96_77 11.551961
Rsn95_77 sn95_77 sn96_77 11.551961
Rsp95_78 sp95_78 sp96_78 11.551961
Rsn95_78 sn95_78 sn96_78 11.551961
Rsp95_79 sp95_79 sp96_79 11.551961
Rsn95_79 sn95_79 sn96_79 11.551961
Rsp95_80 sp95_80 sp96_80 11.551961
Rsn95_80 sn95_80 sn96_80 11.551961
Rsp95_81 sp95_81 sp96_81 11.551961
Rsn95_81 sn95_81 sn96_81 11.551961
Rsp95_82 sp95_82 sp96_82 11.551961
Rsn95_82 sn95_82 sn96_82 11.551961
Rsp95_83 sp95_83 sp96_83 11.551961
Rsn95_83 sn95_83 sn96_83 11.551961
Rsp95_84 sp95_84 sp96_84 11.551961
Rsn95_84 sn95_84 sn96_84 11.551961
Rsp96_1 sp96_1 sp97_1 11.551961
Rsn96_1 sn96_1 sn97_1 11.551961
Rsp96_2 sp96_2 sp97_2 11.551961
Rsn96_2 sn96_2 sn97_2 11.551961
Rsp96_3 sp96_3 sp97_3 11.551961
Rsn96_3 sn96_3 sn97_3 11.551961
Rsp96_4 sp96_4 sp97_4 11.551961
Rsn96_4 sn96_4 sn97_4 11.551961
Rsp96_5 sp96_5 sp97_5 11.551961
Rsn96_5 sn96_5 sn97_5 11.551961
Rsp96_6 sp96_6 sp97_6 11.551961
Rsn96_6 sn96_6 sn97_6 11.551961
Rsp96_7 sp96_7 sp97_7 11.551961
Rsn96_7 sn96_7 sn97_7 11.551961
Rsp96_8 sp96_8 sp97_8 11.551961
Rsn96_8 sn96_8 sn97_8 11.551961
Rsp96_9 sp96_9 sp97_9 11.551961
Rsn96_9 sn96_9 sn97_9 11.551961
Rsp96_10 sp96_10 sp97_10 11.551961
Rsn96_10 sn96_10 sn97_10 11.551961
Rsp96_11 sp96_11 sp97_11 11.551961
Rsn96_11 sn96_11 sn97_11 11.551961
Rsp96_12 sp96_12 sp97_12 11.551961
Rsn96_12 sn96_12 sn97_12 11.551961
Rsp96_13 sp96_13 sp97_13 11.551961
Rsn96_13 sn96_13 sn97_13 11.551961
Rsp96_14 sp96_14 sp97_14 11.551961
Rsn96_14 sn96_14 sn97_14 11.551961
Rsp96_15 sp96_15 sp97_15 11.551961
Rsn96_15 sn96_15 sn97_15 11.551961
Rsp96_16 sp96_16 sp97_16 11.551961
Rsn96_16 sn96_16 sn97_16 11.551961
Rsp96_17 sp96_17 sp97_17 11.551961
Rsn96_17 sn96_17 sn97_17 11.551961
Rsp96_18 sp96_18 sp97_18 11.551961
Rsn96_18 sn96_18 sn97_18 11.551961
Rsp96_19 sp96_19 sp97_19 11.551961
Rsn96_19 sn96_19 sn97_19 11.551961
Rsp96_20 sp96_20 sp97_20 11.551961
Rsn96_20 sn96_20 sn97_20 11.551961
Rsp96_21 sp96_21 sp97_21 11.551961
Rsn96_21 sn96_21 sn97_21 11.551961
Rsp96_22 sp96_22 sp97_22 11.551961
Rsn96_22 sn96_22 sn97_22 11.551961
Rsp96_23 sp96_23 sp97_23 11.551961
Rsn96_23 sn96_23 sn97_23 11.551961
Rsp96_24 sp96_24 sp97_24 11.551961
Rsn96_24 sn96_24 sn97_24 11.551961
Rsp96_25 sp96_25 sp97_25 11.551961
Rsn96_25 sn96_25 sn97_25 11.551961
Rsp96_26 sp96_26 sp97_26 11.551961
Rsn96_26 sn96_26 sn97_26 11.551961
Rsp96_27 sp96_27 sp97_27 11.551961
Rsn96_27 sn96_27 sn97_27 11.551961
Rsp96_28 sp96_28 sp97_28 11.551961
Rsn96_28 sn96_28 sn97_28 11.551961
Rsp96_29 sp96_29 sp97_29 11.551961
Rsn96_29 sn96_29 sn97_29 11.551961
Rsp96_30 sp96_30 sp97_30 11.551961
Rsn96_30 sn96_30 sn97_30 11.551961
Rsp96_31 sp96_31 sp97_31 11.551961
Rsn96_31 sn96_31 sn97_31 11.551961
Rsp96_32 sp96_32 sp97_32 11.551961
Rsn96_32 sn96_32 sn97_32 11.551961
Rsp96_33 sp96_33 sp97_33 11.551961
Rsn96_33 sn96_33 sn97_33 11.551961
Rsp96_34 sp96_34 sp97_34 11.551961
Rsn96_34 sn96_34 sn97_34 11.551961
Rsp96_35 sp96_35 sp97_35 11.551961
Rsn96_35 sn96_35 sn97_35 11.551961
Rsp96_36 sp96_36 sp97_36 11.551961
Rsn96_36 sn96_36 sn97_36 11.551961
Rsp96_37 sp96_37 sp97_37 11.551961
Rsn96_37 sn96_37 sn97_37 11.551961
Rsp96_38 sp96_38 sp97_38 11.551961
Rsn96_38 sn96_38 sn97_38 11.551961
Rsp96_39 sp96_39 sp97_39 11.551961
Rsn96_39 sn96_39 sn97_39 11.551961
Rsp96_40 sp96_40 sp97_40 11.551961
Rsn96_40 sn96_40 sn97_40 11.551961
Rsp96_41 sp96_41 sp97_41 11.551961
Rsn96_41 sn96_41 sn97_41 11.551961
Rsp96_42 sp96_42 sp97_42 11.551961
Rsn96_42 sn96_42 sn97_42 11.551961
Rsp96_43 sp96_43 sp97_43 11.551961
Rsn96_43 sn96_43 sn97_43 11.551961
Rsp96_44 sp96_44 sp97_44 11.551961
Rsn96_44 sn96_44 sn97_44 11.551961
Rsp96_45 sp96_45 sp97_45 11.551961
Rsn96_45 sn96_45 sn97_45 11.551961
Rsp96_46 sp96_46 sp97_46 11.551961
Rsn96_46 sn96_46 sn97_46 11.551961
Rsp96_47 sp96_47 sp97_47 11.551961
Rsn96_47 sn96_47 sn97_47 11.551961
Rsp96_48 sp96_48 sp97_48 11.551961
Rsn96_48 sn96_48 sn97_48 11.551961
Rsp96_49 sp96_49 sp97_49 11.551961
Rsn96_49 sn96_49 sn97_49 11.551961
Rsp96_50 sp96_50 sp97_50 11.551961
Rsn96_50 sn96_50 sn97_50 11.551961
Rsp96_51 sp96_51 sp97_51 11.551961
Rsn96_51 sn96_51 sn97_51 11.551961
Rsp96_52 sp96_52 sp97_52 11.551961
Rsn96_52 sn96_52 sn97_52 11.551961
Rsp96_53 sp96_53 sp97_53 11.551961
Rsn96_53 sn96_53 sn97_53 11.551961
Rsp96_54 sp96_54 sp97_54 11.551961
Rsn96_54 sn96_54 sn97_54 11.551961
Rsp96_55 sp96_55 sp97_55 11.551961
Rsn96_55 sn96_55 sn97_55 11.551961
Rsp96_56 sp96_56 sp97_56 11.551961
Rsn96_56 sn96_56 sn97_56 11.551961
Rsp96_57 sp96_57 sp97_57 11.551961
Rsn96_57 sn96_57 sn97_57 11.551961
Rsp96_58 sp96_58 sp97_58 11.551961
Rsn96_58 sn96_58 sn97_58 11.551961
Rsp96_59 sp96_59 sp97_59 11.551961
Rsn96_59 sn96_59 sn97_59 11.551961
Rsp96_60 sp96_60 sp97_60 11.551961
Rsn96_60 sn96_60 sn97_60 11.551961
Rsp96_61 sp96_61 sp97_61 11.551961
Rsn96_61 sn96_61 sn97_61 11.551961
Rsp96_62 sp96_62 sp97_62 11.551961
Rsn96_62 sn96_62 sn97_62 11.551961
Rsp96_63 sp96_63 sp97_63 11.551961
Rsn96_63 sn96_63 sn97_63 11.551961
Rsp96_64 sp96_64 sp97_64 11.551961
Rsn96_64 sn96_64 sn97_64 11.551961
Rsp96_65 sp96_65 sp97_65 11.551961
Rsn96_65 sn96_65 sn97_65 11.551961
Rsp96_66 sp96_66 sp97_66 11.551961
Rsn96_66 sn96_66 sn97_66 11.551961
Rsp96_67 sp96_67 sp97_67 11.551961
Rsn96_67 sn96_67 sn97_67 11.551961
Rsp96_68 sp96_68 sp97_68 11.551961
Rsn96_68 sn96_68 sn97_68 11.551961
Rsp96_69 sp96_69 sp97_69 11.551961
Rsn96_69 sn96_69 sn97_69 11.551961
Rsp96_70 sp96_70 sp97_70 11.551961
Rsn96_70 sn96_70 sn97_70 11.551961
Rsp96_71 sp96_71 sp97_71 11.551961
Rsn96_71 sn96_71 sn97_71 11.551961
Rsp96_72 sp96_72 sp97_72 11.551961
Rsn96_72 sn96_72 sn97_72 11.551961
Rsp96_73 sp96_73 sp97_73 11.551961
Rsn96_73 sn96_73 sn97_73 11.551961
Rsp96_74 sp96_74 sp97_74 11.551961
Rsn96_74 sn96_74 sn97_74 11.551961
Rsp96_75 sp96_75 sp97_75 11.551961
Rsn96_75 sn96_75 sn97_75 11.551961
Rsp96_76 sp96_76 sp97_76 11.551961
Rsn96_76 sn96_76 sn97_76 11.551961
Rsp96_77 sp96_77 sp97_77 11.551961
Rsn96_77 sn96_77 sn97_77 11.551961
Rsp96_78 sp96_78 sp97_78 11.551961
Rsn96_78 sn96_78 sn97_78 11.551961
Rsp96_79 sp96_79 sp97_79 11.551961
Rsn96_79 sn96_79 sn97_79 11.551961
Rsp96_80 sp96_80 sp97_80 11.551961
Rsn96_80 sn96_80 sn97_80 11.551961
Rsp96_81 sp96_81 sp97_81 11.551961
Rsn96_81 sn96_81 sn97_81 11.551961
Rsp96_82 sp96_82 sp97_82 11.551961
Rsn96_82 sn96_82 sn97_82 11.551961
Rsp96_83 sp96_83 sp97_83 11.551961
Rsn96_83 sn96_83 sn97_83 11.551961
Rsp96_84 sp96_84 sp97_84 11.551961
Rsn96_84 sn96_84 sn97_84 11.551961
Rsp97_1 sp97_1 sp98_1 11.551961
Rsn97_1 sn97_1 sn98_1 11.551961
Rsp97_2 sp97_2 sp98_2 11.551961
Rsn97_2 sn97_2 sn98_2 11.551961
Rsp97_3 sp97_3 sp98_3 11.551961
Rsn97_3 sn97_3 sn98_3 11.551961
Rsp97_4 sp97_4 sp98_4 11.551961
Rsn97_4 sn97_4 sn98_4 11.551961
Rsp97_5 sp97_5 sp98_5 11.551961
Rsn97_5 sn97_5 sn98_5 11.551961
Rsp97_6 sp97_6 sp98_6 11.551961
Rsn97_6 sn97_6 sn98_6 11.551961
Rsp97_7 sp97_7 sp98_7 11.551961
Rsn97_7 sn97_7 sn98_7 11.551961
Rsp97_8 sp97_8 sp98_8 11.551961
Rsn97_8 sn97_8 sn98_8 11.551961
Rsp97_9 sp97_9 sp98_9 11.551961
Rsn97_9 sn97_9 sn98_9 11.551961
Rsp97_10 sp97_10 sp98_10 11.551961
Rsn97_10 sn97_10 sn98_10 11.551961
Rsp97_11 sp97_11 sp98_11 11.551961
Rsn97_11 sn97_11 sn98_11 11.551961
Rsp97_12 sp97_12 sp98_12 11.551961
Rsn97_12 sn97_12 sn98_12 11.551961
Rsp97_13 sp97_13 sp98_13 11.551961
Rsn97_13 sn97_13 sn98_13 11.551961
Rsp97_14 sp97_14 sp98_14 11.551961
Rsn97_14 sn97_14 sn98_14 11.551961
Rsp97_15 sp97_15 sp98_15 11.551961
Rsn97_15 sn97_15 sn98_15 11.551961
Rsp97_16 sp97_16 sp98_16 11.551961
Rsn97_16 sn97_16 sn98_16 11.551961
Rsp97_17 sp97_17 sp98_17 11.551961
Rsn97_17 sn97_17 sn98_17 11.551961
Rsp97_18 sp97_18 sp98_18 11.551961
Rsn97_18 sn97_18 sn98_18 11.551961
Rsp97_19 sp97_19 sp98_19 11.551961
Rsn97_19 sn97_19 sn98_19 11.551961
Rsp97_20 sp97_20 sp98_20 11.551961
Rsn97_20 sn97_20 sn98_20 11.551961
Rsp97_21 sp97_21 sp98_21 11.551961
Rsn97_21 sn97_21 sn98_21 11.551961
Rsp97_22 sp97_22 sp98_22 11.551961
Rsn97_22 sn97_22 sn98_22 11.551961
Rsp97_23 sp97_23 sp98_23 11.551961
Rsn97_23 sn97_23 sn98_23 11.551961
Rsp97_24 sp97_24 sp98_24 11.551961
Rsn97_24 sn97_24 sn98_24 11.551961
Rsp97_25 sp97_25 sp98_25 11.551961
Rsn97_25 sn97_25 sn98_25 11.551961
Rsp97_26 sp97_26 sp98_26 11.551961
Rsn97_26 sn97_26 sn98_26 11.551961
Rsp97_27 sp97_27 sp98_27 11.551961
Rsn97_27 sn97_27 sn98_27 11.551961
Rsp97_28 sp97_28 sp98_28 11.551961
Rsn97_28 sn97_28 sn98_28 11.551961
Rsp97_29 sp97_29 sp98_29 11.551961
Rsn97_29 sn97_29 sn98_29 11.551961
Rsp97_30 sp97_30 sp98_30 11.551961
Rsn97_30 sn97_30 sn98_30 11.551961
Rsp97_31 sp97_31 sp98_31 11.551961
Rsn97_31 sn97_31 sn98_31 11.551961
Rsp97_32 sp97_32 sp98_32 11.551961
Rsn97_32 sn97_32 sn98_32 11.551961
Rsp97_33 sp97_33 sp98_33 11.551961
Rsn97_33 sn97_33 sn98_33 11.551961
Rsp97_34 sp97_34 sp98_34 11.551961
Rsn97_34 sn97_34 sn98_34 11.551961
Rsp97_35 sp97_35 sp98_35 11.551961
Rsn97_35 sn97_35 sn98_35 11.551961
Rsp97_36 sp97_36 sp98_36 11.551961
Rsn97_36 sn97_36 sn98_36 11.551961
Rsp97_37 sp97_37 sp98_37 11.551961
Rsn97_37 sn97_37 sn98_37 11.551961
Rsp97_38 sp97_38 sp98_38 11.551961
Rsn97_38 sn97_38 sn98_38 11.551961
Rsp97_39 sp97_39 sp98_39 11.551961
Rsn97_39 sn97_39 sn98_39 11.551961
Rsp97_40 sp97_40 sp98_40 11.551961
Rsn97_40 sn97_40 sn98_40 11.551961
Rsp97_41 sp97_41 sp98_41 11.551961
Rsn97_41 sn97_41 sn98_41 11.551961
Rsp97_42 sp97_42 sp98_42 11.551961
Rsn97_42 sn97_42 sn98_42 11.551961
Rsp97_43 sp97_43 sp98_43 11.551961
Rsn97_43 sn97_43 sn98_43 11.551961
Rsp97_44 sp97_44 sp98_44 11.551961
Rsn97_44 sn97_44 sn98_44 11.551961
Rsp97_45 sp97_45 sp98_45 11.551961
Rsn97_45 sn97_45 sn98_45 11.551961
Rsp97_46 sp97_46 sp98_46 11.551961
Rsn97_46 sn97_46 sn98_46 11.551961
Rsp97_47 sp97_47 sp98_47 11.551961
Rsn97_47 sn97_47 sn98_47 11.551961
Rsp97_48 sp97_48 sp98_48 11.551961
Rsn97_48 sn97_48 sn98_48 11.551961
Rsp97_49 sp97_49 sp98_49 11.551961
Rsn97_49 sn97_49 sn98_49 11.551961
Rsp97_50 sp97_50 sp98_50 11.551961
Rsn97_50 sn97_50 sn98_50 11.551961
Rsp97_51 sp97_51 sp98_51 11.551961
Rsn97_51 sn97_51 sn98_51 11.551961
Rsp97_52 sp97_52 sp98_52 11.551961
Rsn97_52 sn97_52 sn98_52 11.551961
Rsp97_53 sp97_53 sp98_53 11.551961
Rsn97_53 sn97_53 sn98_53 11.551961
Rsp97_54 sp97_54 sp98_54 11.551961
Rsn97_54 sn97_54 sn98_54 11.551961
Rsp97_55 sp97_55 sp98_55 11.551961
Rsn97_55 sn97_55 sn98_55 11.551961
Rsp97_56 sp97_56 sp98_56 11.551961
Rsn97_56 sn97_56 sn98_56 11.551961
Rsp97_57 sp97_57 sp98_57 11.551961
Rsn97_57 sn97_57 sn98_57 11.551961
Rsp97_58 sp97_58 sp98_58 11.551961
Rsn97_58 sn97_58 sn98_58 11.551961
Rsp97_59 sp97_59 sp98_59 11.551961
Rsn97_59 sn97_59 sn98_59 11.551961
Rsp97_60 sp97_60 sp98_60 11.551961
Rsn97_60 sn97_60 sn98_60 11.551961
Rsp97_61 sp97_61 sp98_61 11.551961
Rsn97_61 sn97_61 sn98_61 11.551961
Rsp97_62 sp97_62 sp98_62 11.551961
Rsn97_62 sn97_62 sn98_62 11.551961
Rsp97_63 sp97_63 sp98_63 11.551961
Rsn97_63 sn97_63 sn98_63 11.551961
Rsp97_64 sp97_64 sp98_64 11.551961
Rsn97_64 sn97_64 sn98_64 11.551961
Rsp97_65 sp97_65 sp98_65 11.551961
Rsn97_65 sn97_65 sn98_65 11.551961
Rsp97_66 sp97_66 sp98_66 11.551961
Rsn97_66 sn97_66 sn98_66 11.551961
Rsp97_67 sp97_67 sp98_67 11.551961
Rsn97_67 sn97_67 sn98_67 11.551961
Rsp97_68 sp97_68 sp98_68 11.551961
Rsn97_68 sn97_68 sn98_68 11.551961
Rsp97_69 sp97_69 sp98_69 11.551961
Rsn97_69 sn97_69 sn98_69 11.551961
Rsp97_70 sp97_70 sp98_70 11.551961
Rsn97_70 sn97_70 sn98_70 11.551961
Rsp97_71 sp97_71 sp98_71 11.551961
Rsn97_71 sn97_71 sn98_71 11.551961
Rsp97_72 sp97_72 sp98_72 11.551961
Rsn97_72 sn97_72 sn98_72 11.551961
Rsp97_73 sp97_73 sp98_73 11.551961
Rsn97_73 sn97_73 sn98_73 11.551961
Rsp97_74 sp97_74 sp98_74 11.551961
Rsn97_74 sn97_74 sn98_74 11.551961
Rsp97_75 sp97_75 sp98_75 11.551961
Rsn97_75 sn97_75 sn98_75 11.551961
Rsp97_76 sp97_76 sp98_76 11.551961
Rsn97_76 sn97_76 sn98_76 11.551961
Rsp97_77 sp97_77 sp98_77 11.551961
Rsn97_77 sn97_77 sn98_77 11.551961
Rsp97_78 sp97_78 sp98_78 11.551961
Rsn97_78 sn97_78 sn98_78 11.551961
Rsp97_79 sp97_79 sp98_79 11.551961
Rsn97_79 sn97_79 sn98_79 11.551961
Rsp97_80 sp97_80 sp98_80 11.551961
Rsn97_80 sn97_80 sn98_80 11.551961
Rsp97_81 sp97_81 sp98_81 11.551961
Rsn97_81 sn97_81 sn98_81 11.551961
Rsp97_82 sp97_82 sp98_82 11.551961
Rsn97_82 sn97_82 sn98_82 11.551961
Rsp97_83 sp97_83 sp98_83 11.551961
Rsn97_83 sn97_83 sn98_83 11.551961
Rsp97_84 sp97_84 sp98_84 11.551961
Rsn97_84 sn97_84 sn98_84 11.551961
Rsp98_1 sp98_1 sp99_1 11.551961
Rsn98_1 sn98_1 sn99_1 11.551961
Rsp98_2 sp98_2 sp99_2 11.551961
Rsn98_2 sn98_2 sn99_2 11.551961
Rsp98_3 sp98_3 sp99_3 11.551961
Rsn98_3 sn98_3 sn99_3 11.551961
Rsp98_4 sp98_4 sp99_4 11.551961
Rsn98_4 sn98_4 sn99_4 11.551961
Rsp98_5 sp98_5 sp99_5 11.551961
Rsn98_5 sn98_5 sn99_5 11.551961
Rsp98_6 sp98_6 sp99_6 11.551961
Rsn98_6 sn98_6 sn99_6 11.551961
Rsp98_7 sp98_7 sp99_7 11.551961
Rsn98_7 sn98_7 sn99_7 11.551961
Rsp98_8 sp98_8 sp99_8 11.551961
Rsn98_8 sn98_8 sn99_8 11.551961
Rsp98_9 sp98_9 sp99_9 11.551961
Rsn98_9 sn98_9 sn99_9 11.551961
Rsp98_10 sp98_10 sp99_10 11.551961
Rsn98_10 sn98_10 sn99_10 11.551961
Rsp98_11 sp98_11 sp99_11 11.551961
Rsn98_11 sn98_11 sn99_11 11.551961
Rsp98_12 sp98_12 sp99_12 11.551961
Rsn98_12 sn98_12 sn99_12 11.551961
Rsp98_13 sp98_13 sp99_13 11.551961
Rsn98_13 sn98_13 sn99_13 11.551961
Rsp98_14 sp98_14 sp99_14 11.551961
Rsn98_14 sn98_14 sn99_14 11.551961
Rsp98_15 sp98_15 sp99_15 11.551961
Rsn98_15 sn98_15 sn99_15 11.551961
Rsp98_16 sp98_16 sp99_16 11.551961
Rsn98_16 sn98_16 sn99_16 11.551961
Rsp98_17 sp98_17 sp99_17 11.551961
Rsn98_17 sn98_17 sn99_17 11.551961
Rsp98_18 sp98_18 sp99_18 11.551961
Rsn98_18 sn98_18 sn99_18 11.551961
Rsp98_19 sp98_19 sp99_19 11.551961
Rsn98_19 sn98_19 sn99_19 11.551961
Rsp98_20 sp98_20 sp99_20 11.551961
Rsn98_20 sn98_20 sn99_20 11.551961
Rsp98_21 sp98_21 sp99_21 11.551961
Rsn98_21 sn98_21 sn99_21 11.551961
Rsp98_22 sp98_22 sp99_22 11.551961
Rsn98_22 sn98_22 sn99_22 11.551961
Rsp98_23 sp98_23 sp99_23 11.551961
Rsn98_23 sn98_23 sn99_23 11.551961
Rsp98_24 sp98_24 sp99_24 11.551961
Rsn98_24 sn98_24 sn99_24 11.551961
Rsp98_25 sp98_25 sp99_25 11.551961
Rsn98_25 sn98_25 sn99_25 11.551961
Rsp98_26 sp98_26 sp99_26 11.551961
Rsn98_26 sn98_26 sn99_26 11.551961
Rsp98_27 sp98_27 sp99_27 11.551961
Rsn98_27 sn98_27 sn99_27 11.551961
Rsp98_28 sp98_28 sp99_28 11.551961
Rsn98_28 sn98_28 sn99_28 11.551961
Rsp98_29 sp98_29 sp99_29 11.551961
Rsn98_29 sn98_29 sn99_29 11.551961
Rsp98_30 sp98_30 sp99_30 11.551961
Rsn98_30 sn98_30 sn99_30 11.551961
Rsp98_31 sp98_31 sp99_31 11.551961
Rsn98_31 sn98_31 sn99_31 11.551961
Rsp98_32 sp98_32 sp99_32 11.551961
Rsn98_32 sn98_32 sn99_32 11.551961
Rsp98_33 sp98_33 sp99_33 11.551961
Rsn98_33 sn98_33 sn99_33 11.551961
Rsp98_34 sp98_34 sp99_34 11.551961
Rsn98_34 sn98_34 sn99_34 11.551961
Rsp98_35 sp98_35 sp99_35 11.551961
Rsn98_35 sn98_35 sn99_35 11.551961
Rsp98_36 sp98_36 sp99_36 11.551961
Rsn98_36 sn98_36 sn99_36 11.551961
Rsp98_37 sp98_37 sp99_37 11.551961
Rsn98_37 sn98_37 sn99_37 11.551961
Rsp98_38 sp98_38 sp99_38 11.551961
Rsn98_38 sn98_38 sn99_38 11.551961
Rsp98_39 sp98_39 sp99_39 11.551961
Rsn98_39 sn98_39 sn99_39 11.551961
Rsp98_40 sp98_40 sp99_40 11.551961
Rsn98_40 sn98_40 sn99_40 11.551961
Rsp98_41 sp98_41 sp99_41 11.551961
Rsn98_41 sn98_41 sn99_41 11.551961
Rsp98_42 sp98_42 sp99_42 11.551961
Rsn98_42 sn98_42 sn99_42 11.551961
Rsp98_43 sp98_43 sp99_43 11.551961
Rsn98_43 sn98_43 sn99_43 11.551961
Rsp98_44 sp98_44 sp99_44 11.551961
Rsn98_44 sn98_44 sn99_44 11.551961
Rsp98_45 sp98_45 sp99_45 11.551961
Rsn98_45 sn98_45 sn99_45 11.551961
Rsp98_46 sp98_46 sp99_46 11.551961
Rsn98_46 sn98_46 sn99_46 11.551961
Rsp98_47 sp98_47 sp99_47 11.551961
Rsn98_47 sn98_47 sn99_47 11.551961
Rsp98_48 sp98_48 sp99_48 11.551961
Rsn98_48 sn98_48 sn99_48 11.551961
Rsp98_49 sp98_49 sp99_49 11.551961
Rsn98_49 sn98_49 sn99_49 11.551961
Rsp98_50 sp98_50 sp99_50 11.551961
Rsn98_50 sn98_50 sn99_50 11.551961
Rsp98_51 sp98_51 sp99_51 11.551961
Rsn98_51 sn98_51 sn99_51 11.551961
Rsp98_52 sp98_52 sp99_52 11.551961
Rsn98_52 sn98_52 sn99_52 11.551961
Rsp98_53 sp98_53 sp99_53 11.551961
Rsn98_53 sn98_53 sn99_53 11.551961
Rsp98_54 sp98_54 sp99_54 11.551961
Rsn98_54 sn98_54 sn99_54 11.551961
Rsp98_55 sp98_55 sp99_55 11.551961
Rsn98_55 sn98_55 sn99_55 11.551961
Rsp98_56 sp98_56 sp99_56 11.551961
Rsn98_56 sn98_56 sn99_56 11.551961
Rsp98_57 sp98_57 sp99_57 11.551961
Rsn98_57 sn98_57 sn99_57 11.551961
Rsp98_58 sp98_58 sp99_58 11.551961
Rsn98_58 sn98_58 sn99_58 11.551961
Rsp98_59 sp98_59 sp99_59 11.551961
Rsn98_59 sn98_59 sn99_59 11.551961
Rsp98_60 sp98_60 sp99_60 11.551961
Rsn98_60 sn98_60 sn99_60 11.551961
Rsp98_61 sp98_61 sp99_61 11.551961
Rsn98_61 sn98_61 sn99_61 11.551961
Rsp98_62 sp98_62 sp99_62 11.551961
Rsn98_62 sn98_62 sn99_62 11.551961
Rsp98_63 sp98_63 sp99_63 11.551961
Rsn98_63 sn98_63 sn99_63 11.551961
Rsp98_64 sp98_64 sp99_64 11.551961
Rsn98_64 sn98_64 sn99_64 11.551961
Rsp98_65 sp98_65 sp99_65 11.551961
Rsn98_65 sn98_65 sn99_65 11.551961
Rsp98_66 sp98_66 sp99_66 11.551961
Rsn98_66 sn98_66 sn99_66 11.551961
Rsp98_67 sp98_67 sp99_67 11.551961
Rsn98_67 sn98_67 sn99_67 11.551961
Rsp98_68 sp98_68 sp99_68 11.551961
Rsn98_68 sn98_68 sn99_68 11.551961
Rsp98_69 sp98_69 sp99_69 11.551961
Rsn98_69 sn98_69 sn99_69 11.551961
Rsp98_70 sp98_70 sp99_70 11.551961
Rsn98_70 sn98_70 sn99_70 11.551961
Rsp98_71 sp98_71 sp99_71 11.551961
Rsn98_71 sn98_71 sn99_71 11.551961
Rsp98_72 sp98_72 sp99_72 11.551961
Rsn98_72 sn98_72 sn99_72 11.551961
Rsp98_73 sp98_73 sp99_73 11.551961
Rsn98_73 sn98_73 sn99_73 11.551961
Rsp98_74 sp98_74 sp99_74 11.551961
Rsn98_74 sn98_74 sn99_74 11.551961
Rsp98_75 sp98_75 sp99_75 11.551961
Rsn98_75 sn98_75 sn99_75 11.551961
Rsp98_76 sp98_76 sp99_76 11.551961
Rsn98_76 sn98_76 sn99_76 11.551961
Rsp98_77 sp98_77 sp99_77 11.551961
Rsn98_77 sn98_77 sn99_77 11.551961
Rsp98_78 sp98_78 sp99_78 11.551961
Rsn98_78 sn98_78 sn99_78 11.551961
Rsp98_79 sp98_79 sp99_79 11.551961
Rsn98_79 sn98_79 sn99_79 11.551961
Rsp98_80 sp98_80 sp99_80 11.551961
Rsn98_80 sn98_80 sn99_80 11.551961
Rsp98_81 sp98_81 sp99_81 11.551961
Rsn98_81 sn98_81 sn99_81 11.551961
Rsp98_82 sp98_82 sp99_82 11.551961
Rsn98_82 sn98_82 sn99_82 11.551961
Rsp98_83 sp98_83 sp99_83 11.551961
Rsn98_83 sn98_83 sn99_83 11.551961
Rsp98_84 sp98_84 sp99_84 11.551961
Rsn98_84 sn98_84 sn99_84 11.551961
Rsp99_1 sp99_1 sp100_1 11.551961
Rsn99_1 sn99_1 sn100_1 11.551961
Rsp99_2 sp99_2 sp100_2 11.551961
Rsn99_2 sn99_2 sn100_2 11.551961
Rsp99_3 sp99_3 sp100_3 11.551961
Rsn99_3 sn99_3 sn100_3 11.551961
Rsp99_4 sp99_4 sp100_4 11.551961
Rsn99_4 sn99_4 sn100_4 11.551961
Rsp99_5 sp99_5 sp100_5 11.551961
Rsn99_5 sn99_5 sn100_5 11.551961
Rsp99_6 sp99_6 sp100_6 11.551961
Rsn99_6 sn99_6 sn100_6 11.551961
Rsp99_7 sp99_7 sp100_7 11.551961
Rsn99_7 sn99_7 sn100_7 11.551961
Rsp99_8 sp99_8 sp100_8 11.551961
Rsn99_8 sn99_8 sn100_8 11.551961
Rsp99_9 sp99_9 sp100_9 11.551961
Rsn99_9 sn99_9 sn100_9 11.551961
Rsp99_10 sp99_10 sp100_10 11.551961
Rsn99_10 sn99_10 sn100_10 11.551961
Rsp99_11 sp99_11 sp100_11 11.551961
Rsn99_11 sn99_11 sn100_11 11.551961
Rsp99_12 sp99_12 sp100_12 11.551961
Rsn99_12 sn99_12 sn100_12 11.551961
Rsp99_13 sp99_13 sp100_13 11.551961
Rsn99_13 sn99_13 sn100_13 11.551961
Rsp99_14 sp99_14 sp100_14 11.551961
Rsn99_14 sn99_14 sn100_14 11.551961
Rsp99_15 sp99_15 sp100_15 11.551961
Rsn99_15 sn99_15 sn100_15 11.551961
Rsp99_16 sp99_16 sp100_16 11.551961
Rsn99_16 sn99_16 sn100_16 11.551961
Rsp99_17 sp99_17 sp100_17 11.551961
Rsn99_17 sn99_17 sn100_17 11.551961
Rsp99_18 sp99_18 sp100_18 11.551961
Rsn99_18 sn99_18 sn100_18 11.551961
Rsp99_19 sp99_19 sp100_19 11.551961
Rsn99_19 sn99_19 sn100_19 11.551961
Rsp99_20 sp99_20 sp100_20 11.551961
Rsn99_20 sn99_20 sn100_20 11.551961
Rsp99_21 sp99_21 sp100_21 11.551961
Rsn99_21 sn99_21 sn100_21 11.551961
Rsp99_22 sp99_22 sp100_22 11.551961
Rsn99_22 sn99_22 sn100_22 11.551961
Rsp99_23 sp99_23 sp100_23 11.551961
Rsn99_23 sn99_23 sn100_23 11.551961
Rsp99_24 sp99_24 sp100_24 11.551961
Rsn99_24 sn99_24 sn100_24 11.551961
Rsp99_25 sp99_25 sp100_25 11.551961
Rsn99_25 sn99_25 sn100_25 11.551961
Rsp99_26 sp99_26 sp100_26 11.551961
Rsn99_26 sn99_26 sn100_26 11.551961
Rsp99_27 sp99_27 sp100_27 11.551961
Rsn99_27 sn99_27 sn100_27 11.551961
Rsp99_28 sp99_28 sp100_28 11.551961
Rsn99_28 sn99_28 sn100_28 11.551961
Rsp99_29 sp99_29 sp100_29 11.551961
Rsn99_29 sn99_29 sn100_29 11.551961
Rsp99_30 sp99_30 sp100_30 11.551961
Rsn99_30 sn99_30 sn100_30 11.551961
Rsp99_31 sp99_31 sp100_31 11.551961
Rsn99_31 sn99_31 sn100_31 11.551961
Rsp99_32 sp99_32 sp100_32 11.551961
Rsn99_32 sn99_32 sn100_32 11.551961
Rsp99_33 sp99_33 sp100_33 11.551961
Rsn99_33 sn99_33 sn100_33 11.551961
Rsp99_34 sp99_34 sp100_34 11.551961
Rsn99_34 sn99_34 sn100_34 11.551961
Rsp99_35 sp99_35 sp100_35 11.551961
Rsn99_35 sn99_35 sn100_35 11.551961
Rsp99_36 sp99_36 sp100_36 11.551961
Rsn99_36 sn99_36 sn100_36 11.551961
Rsp99_37 sp99_37 sp100_37 11.551961
Rsn99_37 sn99_37 sn100_37 11.551961
Rsp99_38 sp99_38 sp100_38 11.551961
Rsn99_38 sn99_38 sn100_38 11.551961
Rsp99_39 sp99_39 sp100_39 11.551961
Rsn99_39 sn99_39 sn100_39 11.551961
Rsp99_40 sp99_40 sp100_40 11.551961
Rsn99_40 sn99_40 sn100_40 11.551961
Rsp99_41 sp99_41 sp100_41 11.551961
Rsn99_41 sn99_41 sn100_41 11.551961
Rsp99_42 sp99_42 sp100_42 11.551961
Rsn99_42 sn99_42 sn100_42 11.551961
Rsp99_43 sp99_43 sp100_43 11.551961
Rsn99_43 sn99_43 sn100_43 11.551961
Rsp99_44 sp99_44 sp100_44 11.551961
Rsn99_44 sn99_44 sn100_44 11.551961
Rsp99_45 sp99_45 sp100_45 11.551961
Rsn99_45 sn99_45 sn100_45 11.551961
Rsp99_46 sp99_46 sp100_46 11.551961
Rsn99_46 sn99_46 sn100_46 11.551961
Rsp99_47 sp99_47 sp100_47 11.551961
Rsn99_47 sn99_47 sn100_47 11.551961
Rsp99_48 sp99_48 sp100_48 11.551961
Rsn99_48 sn99_48 sn100_48 11.551961
Rsp99_49 sp99_49 sp100_49 11.551961
Rsn99_49 sn99_49 sn100_49 11.551961
Rsp99_50 sp99_50 sp100_50 11.551961
Rsn99_50 sn99_50 sn100_50 11.551961
Rsp99_51 sp99_51 sp100_51 11.551961
Rsn99_51 sn99_51 sn100_51 11.551961
Rsp99_52 sp99_52 sp100_52 11.551961
Rsn99_52 sn99_52 sn100_52 11.551961
Rsp99_53 sp99_53 sp100_53 11.551961
Rsn99_53 sn99_53 sn100_53 11.551961
Rsp99_54 sp99_54 sp100_54 11.551961
Rsn99_54 sn99_54 sn100_54 11.551961
Rsp99_55 sp99_55 sp100_55 11.551961
Rsn99_55 sn99_55 sn100_55 11.551961
Rsp99_56 sp99_56 sp100_56 11.551961
Rsn99_56 sn99_56 sn100_56 11.551961
Rsp99_57 sp99_57 sp100_57 11.551961
Rsn99_57 sn99_57 sn100_57 11.551961
Rsp99_58 sp99_58 sp100_58 11.551961
Rsn99_58 sn99_58 sn100_58 11.551961
Rsp99_59 sp99_59 sp100_59 11.551961
Rsn99_59 sn99_59 sn100_59 11.551961
Rsp99_60 sp99_60 sp100_60 11.551961
Rsn99_60 sn99_60 sn100_60 11.551961
Rsp99_61 sp99_61 sp100_61 11.551961
Rsn99_61 sn99_61 sn100_61 11.551961
Rsp99_62 sp99_62 sp100_62 11.551961
Rsn99_62 sn99_62 sn100_62 11.551961
Rsp99_63 sp99_63 sp100_63 11.551961
Rsn99_63 sn99_63 sn100_63 11.551961
Rsp99_64 sp99_64 sp100_64 11.551961
Rsn99_64 sn99_64 sn100_64 11.551961
Rsp99_65 sp99_65 sp100_65 11.551961
Rsn99_65 sn99_65 sn100_65 11.551961
Rsp99_66 sp99_66 sp100_66 11.551961
Rsn99_66 sn99_66 sn100_66 11.551961
Rsp99_67 sp99_67 sp100_67 11.551961
Rsn99_67 sn99_67 sn100_67 11.551961
Rsp99_68 sp99_68 sp100_68 11.551961
Rsn99_68 sn99_68 sn100_68 11.551961
Rsp99_69 sp99_69 sp100_69 11.551961
Rsn99_69 sn99_69 sn100_69 11.551961
Rsp99_70 sp99_70 sp100_70 11.551961
Rsn99_70 sn99_70 sn100_70 11.551961
Rsp99_71 sp99_71 sp100_71 11.551961
Rsn99_71 sn99_71 sn100_71 11.551961
Rsp99_72 sp99_72 sp100_72 11.551961
Rsn99_72 sn99_72 sn100_72 11.551961
Rsp99_73 sp99_73 sp100_73 11.551961
Rsn99_73 sn99_73 sn100_73 11.551961
Rsp99_74 sp99_74 sp100_74 11.551961
Rsn99_74 sn99_74 sn100_74 11.551961
Rsp99_75 sp99_75 sp100_75 11.551961
Rsn99_75 sn99_75 sn100_75 11.551961
Rsp99_76 sp99_76 sp100_76 11.551961
Rsn99_76 sn99_76 sn100_76 11.551961
Rsp99_77 sp99_77 sp100_77 11.551961
Rsn99_77 sn99_77 sn100_77 11.551961
Rsp99_78 sp99_78 sp100_78 11.551961
Rsn99_78 sn99_78 sn100_78 11.551961
Rsp99_79 sp99_79 sp100_79 11.551961
Rsn99_79 sn99_79 sn100_79 11.551961
Rsp99_80 sp99_80 sp100_80 11.551961
Rsn99_80 sn99_80 sn100_80 11.551961
Rsp99_81 sp99_81 sp100_81 11.551961
Rsn99_81 sn99_81 sn100_81 11.551961
Rsp99_82 sp99_82 sp100_82 11.551961
Rsn99_82 sn99_82 sn100_82 11.551961
Rsp99_83 sp99_83 sp100_83 11.551961
Rsn99_83 sn99_83 sn100_83 11.551961
Rsp99_84 sp99_84 sp100_84 11.551961
Rsn99_84 sn99_84 sn100_84 11.551961
Rsp100_1 sp100_1 sp101_1 11.551961
Rsn100_1 sn100_1 sn101_1 11.551961
Rsp100_2 sp100_2 sp101_2 11.551961
Rsn100_2 sn100_2 sn101_2 11.551961
Rsp100_3 sp100_3 sp101_3 11.551961
Rsn100_3 sn100_3 sn101_3 11.551961
Rsp100_4 sp100_4 sp101_4 11.551961
Rsn100_4 sn100_4 sn101_4 11.551961
Rsp100_5 sp100_5 sp101_5 11.551961
Rsn100_5 sn100_5 sn101_5 11.551961
Rsp100_6 sp100_6 sp101_6 11.551961
Rsn100_6 sn100_6 sn101_6 11.551961
Rsp100_7 sp100_7 sp101_7 11.551961
Rsn100_7 sn100_7 sn101_7 11.551961
Rsp100_8 sp100_8 sp101_8 11.551961
Rsn100_8 sn100_8 sn101_8 11.551961
Rsp100_9 sp100_9 sp101_9 11.551961
Rsn100_9 sn100_9 sn101_9 11.551961
Rsp100_10 sp100_10 sp101_10 11.551961
Rsn100_10 sn100_10 sn101_10 11.551961
Rsp100_11 sp100_11 sp101_11 11.551961
Rsn100_11 sn100_11 sn101_11 11.551961
Rsp100_12 sp100_12 sp101_12 11.551961
Rsn100_12 sn100_12 sn101_12 11.551961
Rsp100_13 sp100_13 sp101_13 11.551961
Rsn100_13 sn100_13 sn101_13 11.551961
Rsp100_14 sp100_14 sp101_14 11.551961
Rsn100_14 sn100_14 sn101_14 11.551961
Rsp100_15 sp100_15 sp101_15 11.551961
Rsn100_15 sn100_15 sn101_15 11.551961
Rsp100_16 sp100_16 sp101_16 11.551961
Rsn100_16 sn100_16 sn101_16 11.551961
Rsp100_17 sp100_17 sp101_17 11.551961
Rsn100_17 sn100_17 sn101_17 11.551961
Rsp100_18 sp100_18 sp101_18 11.551961
Rsn100_18 sn100_18 sn101_18 11.551961
Rsp100_19 sp100_19 sp101_19 11.551961
Rsn100_19 sn100_19 sn101_19 11.551961
Rsp100_20 sp100_20 sp101_20 11.551961
Rsn100_20 sn100_20 sn101_20 11.551961
Rsp100_21 sp100_21 sp101_21 11.551961
Rsn100_21 sn100_21 sn101_21 11.551961
Rsp100_22 sp100_22 sp101_22 11.551961
Rsn100_22 sn100_22 sn101_22 11.551961
Rsp100_23 sp100_23 sp101_23 11.551961
Rsn100_23 sn100_23 sn101_23 11.551961
Rsp100_24 sp100_24 sp101_24 11.551961
Rsn100_24 sn100_24 sn101_24 11.551961
Rsp100_25 sp100_25 sp101_25 11.551961
Rsn100_25 sn100_25 sn101_25 11.551961
Rsp100_26 sp100_26 sp101_26 11.551961
Rsn100_26 sn100_26 sn101_26 11.551961
Rsp100_27 sp100_27 sp101_27 11.551961
Rsn100_27 sn100_27 sn101_27 11.551961
Rsp100_28 sp100_28 sp101_28 11.551961
Rsn100_28 sn100_28 sn101_28 11.551961
Rsp100_29 sp100_29 sp101_29 11.551961
Rsn100_29 sn100_29 sn101_29 11.551961
Rsp100_30 sp100_30 sp101_30 11.551961
Rsn100_30 sn100_30 sn101_30 11.551961
Rsp100_31 sp100_31 sp101_31 11.551961
Rsn100_31 sn100_31 sn101_31 11.551961
Rsp100_32 sp100_32 sp101_32 11.551961
Rsn100_32 sn100_32 sn101_32 11.551961
Rsp100_33 sp100_33 sp101_33 11.551961
Rsn100_33 sn100_33 sn101_33 11.551961
Rsp100_34 sp100_34 sp101_34 11.551961
Rsn100_34 sn100_34 sn101_34 11.551961
Rsp100_35 sp100_35 sp101_35 11.551961
Rsn100_35 sn100_35 sn101_35 11.551961
Rsp100_36 sp100_36 sp101_36 11.551961
Rsn100_36 sn100_36 sn101_36 11.551961
Rsp100_37 sp100_37 sp101_37 11.551961
Rsn100_37 sn100_37 sn101_37 11.551961
Rsp100_38 sp100_38 sp101_38 11.551961
Rsn100_38 sn100_38 sn101_38 11.551961
Rsp100_39 sp100_39 sp101_39 11.551961
Rsn100_39 sn100_39 sn101_39 11.551961
Rsp100_40 sp100_40 sp101_40 11.551961
Rsn100_40 sn100_40 sn101_40 11.551961
Rsp100_41 sp100_41 sp101_41 11.551961
Rsn100_41 sn100_41 sn101_41 11.551961
Rsp100_42 sp100_42 sp101_42 11.551961
Rsn100_42 sn100_42 sn101_42 11.551961
Rsp100_43 sp100_43 sp101_43 11.551961
Rsn100_43 sn100_43 sn101_43 11.551961
Rsp100_44 sp100_44 sp101_44 11.551961
Rsn100_44 sn100_44 sn101_44 11.551961
Rsp100_45 sp100_45 sp101_45 11.551961
Rsn100_45 sn100_45 sn101_45 11.551961
Rsp100_46 sp100_46 sp101_46 11.551961
Rsn100_46 sn100_46 sn101_46 11.551961
Rsp100_47 sp100_47 sp101_47 11.551961
Rsn100_47 sn100_47 sn101_47 11.551961
Rsp100_48 sp100_48 sp101_48 11.551961
Rsn100_48 sn100_48 sn101_48 11.551961
Rsp100_49 sp100_49 sp101_49 11.551961
Rsn100_49 sn100_49 sn101_49 11.551961
Rsp100_50 sp100_50 sp101_50 11.551961
Rsn100_50 sn100_50 sn101_50 11.551961
Rsp100_51 sp100_51 sp101_51 11.551961
Rsn100_51 sn100_51 sn101_51 11.551961
Rsp100_52 sp100_52 sp101_52 11.551961
Rsn100_52 sn100_52 sn101_52 11.551961
Rsp100_53 sp100_53 sp101_53 11.551961
Rsn100_53 sn100_53 sn101_53 11.551961
Rsp100_54 sp100_54 sp101_54 11.551961
Rsn100_54 sn100_54 sn101_54 11.551961
Rsp100_55 sp100_55 sp101_55 11.551961
Rsn100_55 sn100_55 sn101_55 11.551961
Rsp100_56 sp100_56 sp101_56 11.551961
Rsn100_56 sn100_56 sn101_56 11.551961
Rsp100_57 sp100_57 sp101_57 11.551961
Rsn100_57 sn100_57 sn101_57 11.551961
Rsp100_58 sp100_58 sp101_58 11.551961
Rsn100_58 sn100_58 sn101_58 11.551961
Rsp100_59 sp100_59 sp101_59 11.551961
Rsn100_59 sn100_59 sn101_59 11.551961
Rsp100_60 sp100_60 sp101_60 11.551961
Rsn100_60 sn100_60 sn101_60 11.551961
Rsp100_61 sp100_61 sp101_61 11.551961
Rsn100_61 sn100_61 sn101_61 11.551961
Rsp100_62 sp100_62 sp101_62 11.551961
Rsn100_62 sn100_62 sn101_62 11.551961
Rsp100_63 sp100_63 sp101_63 11.551961
Rsn100_63 sn100_63 sn101_63 11.551961
Rsp100_64 sp100_64 sp101_64 11.551961
Rsn100_64 sn100_64 sn101_64 11.551961
Rsp100_65 sp100_65 sp101_65 11.551961
Rsn100_65 sn100_65 sn101_65 11.551961
Rsp100_66 sp100_66 sp101_66 11.551961
Rsn100_66 sn100_66 sn101_66 11.551961
Rsp100_67 sp100_67 sp101_67 11.551961
Rsn100_67 sn100_67 sn101_67 11.551961
Rsp100_68 sp100_68 sp101_68 11.551961
Rsn100_68 sn100_68 sn101_68 11.551961
Rsp100_69 sp100_69 sp101_69 11.551961
Rsn100_69 sn100_69 sn101_69 11.551961
Rsp100_70 sp100_70 sp101_70 11.551961
Rsn100_70 sn100_70 sn101_70 11.551961
Rsp100_71 sp100_71 sp101_71 11.551961
Rsn100_71 sn100_71 sn101_71 11.551961
Rsp100_72 sp100_72 sp101_72 11.551961
Rsn100_72 sn100_72 sn101_72 11.551961
Rsp100_73 sp100_73 sp101_73 11.551961
Rsn100_73 sn100_73 sn101_73 11.551961
Rsp100_74 sp100_74 sp101_74 11.551961
Rsn100_74 sn100_74 sn101_74 11.551961
Rsp100_75 sp100_75 sp101_75 11.551961
Rsn100_75 sn100_75 sn101_75 11.551961
Rsp100_76 sp100_76 sp101_76 11.551961
Rsn100_76 sn100_76 sn101_76 11.551961
Rsp100_77 sp100_77 sp101_77 11.551961
Rsn100_77 sn100_77 sn101_77 11.551961
Rsp100_78 sp100_78 sp101_78 11.551961
Rsn100_78 sn100_78 sn101_78 11.551961
Rsp100_79 sp100_79 sp101_79 11.551961
Rsn100_79 sn100_79 sn101_79 11.551961
Rsp100_80 sp100_80 sp101_80 11.551961
Rsn100_80 sn100_80 sn101_80 11.551961
Rsp100_81 sp100_81 sp101_81 11.551961
Rsn100_81 sn100_81 sn101_81 11.551961
Rsp100_82 sp100_82 sp101_82 11.551961
Rsn100_82 sn100_82 sn101_82 11.551961
Rsp100_83 sp100_83 sp101_83 11.551961
Rsn100_83 sn100_83 sn101_83 11.551961
Rsp100_84 sp100_84 sp101_84 11.551961
Rsn100_84 sn100_84 sn101_84 11.551961
Rsp101_1 sp101_1 sp102_1 11.551961
Rsn101_1 sn101_1 sn102_1 11.551961
Rsp101_2 sp101_2 sp102_2 11.551961
Rsn101_2 sn101_2 sn102_2 11.551961
Rsp101_3 sp101_3 sp102_3 11.551961
Rsn101_3 sn101_3 sn102_3 11.551961
Rsp101_4 sp101_4 sp102_4 11.551961
Rsn101_4 sn101_4 sn102_4 11.551961
Rsp101_5 sp101_5 sp102_5 11.551961
Rsn101_5 sn101_5 sn102_5 11.551961
Rsp101_6 sp101_6 sp102_6 11.551961
Rsn101_6 sn101_6 sn102_6 11.551961
Rsp101_7 sp101_7 sp102_7 11.551961
Rsn101_7 sn101_7 sn102_7 11.551961
Rsp101_8 sp101_8 sp102_8 11.551961
Rsn101_8 sn101_8 sn102_8 11.551961
Rsp101_9 sp101_9 sp102_9 11.551961
Rsn101_9 sn101_9 sn102_9 11.551961
Rsp101_10 sp101_10 sp102_10 11.551961
Rsn101_10 sn101_10 sn102_10 11.551961
Rsp101_11 sp101_11 sp102_11 11.551961
Rsn101_11 sn101_11 sn102_11 11.551961
Rsp101_12 sp101_12 sp102_12 11.551961
Rsn101_12 sn101_12 sn102_12 11.551961
Rsp101_13 sp101_13 sp102_13 11.551961
Rsn101_13 sn101_13 sn102_13 11.551961
Rsp101_14 sp101_14 sp102_14 11.551961
Rsn101_14 sn101_14 sn102_14 11.551961
Rsp101_15 sp101_15 sp102_15 11.551961
Rsn101_15 sn101_15 sn102_15 11.551961
Rsp101_16 sp101_16 sp102_16 11.551961
Rsn101_16 sn101_16 sn102_16 11.551961
Rsp101_17 sp101_17 sp102_17 11.551961
Rsn101_17 sn101_17 sn102_17 11.551961
Rsp101_18 sp101_18 sp102_18 11.551961
Rsn101_18 sn101_18 sn102_18 11.551961
Rsp101_19 sp101_19 sp102_19 11.551961
Rsn101_19 sn101_19 sn102_19 11.551961
Rsp101_20 sp101_20 sp102_20 11.551961
Rsn101_20 sn101_20 sn102_20 11.551961
Rsp101_21 sp101_21 sp102_21 11.551961
Rsn101_21 sn101_21 sn102_21 11.551961
Rsp101_22 sp101_22 sp102_22 11.551961
Rsn101_22 sn101_22 sn102_22 11.551961
Rsp101_23 sp101_23 sp102_23 11.551961
Rsn101_23 sn101_23 sn102_23 11.551961
Rsp101_24 sp101_24 sp102_24 11.551961
Rsn101_24 sn101_24 sn102_24 11.551961
Rsp101_25 sp101_25 sp102_25 11.551961
Rsn101_25 sn101_25 sn102_25 11.551961
Rsp101_26 sp101_26 sp102_26 11.551961
Rsn101_26 sn101_26 sn102_26 11.551961
Rsp101_27 sp101_27 sp102_27 11.551961
Rsn101_27 sn101_27 sn102_27 11.551961
Rsp101_28 sp101_28 sp102_28 11.551961
Rsn101_28 sn101_28 sn102_28 11.551961
Rsp101_29 sp101_29 sp102_29 11.551961
Rsn101_29 sn101_29 sn102_29 11.551961
Rsp101_30 sp101_30 sp102_30 11.551961
Rsn101_30 sn101_30 sn102_30 11.551961
Rsp101_31 sp101_31 sp102_31 11.551961
Rsn101_31 sn101_31 sn102_31 11.551961
Rsp101_32 sp101_32 sp102_32 11.551961
Rsn101_32 sn101_32 sn102_32 11.551961
Rsp101_33 sp101_33 sp102_33 11.551961
Rsn101_33 sn101_33 sn102_33 11.551961
Rsp101_34 sp101_34 sp102_34 11.551961
Rsn101_34 sn101_34 sn102_34 11.551961
Rsp101_35 sp101_35 sp102_35 11.551961
Rsn101_35 sn101_35 sn102_35 11.551961
Rsp101_36 sp101_36 sp102_36 11.551961
Rsn101_36 sn101_36 sn102_36 11.551961
Rsp101_37 sp101_37 sp102_37 11.551961
Rsn101_37 sn101_37 sn102_37 11.551961
Rsp101_38 sp101_38 sp102_38 11.551961
Rsn101_38 sn101_38 sn102_38 11.551961
Rsp101_39 sp101_39 sp102_39 11.551961
Rsn101_39 sn101_39 sn102_39 11.551961
Rsp101_40 sp101_40 sp102_40 11.551961
Rsn101_40 sn101_40 sn102_40 11.551961
Rsp101_41 sp101_41 sp102_41 11.551961
Rsn101_41 sn101_41 sn102_41 11.551961
Rsp101_42 sp101_42 sp102_42 11.551961
Rsn101_42 sn101_42 sn102_42 11.551961
Rsp101_43 sp101_43 sp102_43 11.551961
Rsn101_43 sn101_43 sn102_43 11.551961
Rsp101_44 sp101_44 sp102_44 11.551961
Rsn101_44 sn101_44 sn102_44 11.551961
Rsp101_45 sp101_45 sp102_45 11.551961
Rsn101_45 sn101_45 sn102_45 11.551961
Rsp101_46 sp101_46 sp102_46 11.551961
Rsn101_46 sn101_46 sn102_46 11.551961
Rsp101_47 sp101_47 sp102_47 11.551961
Rsn101_47 sn101_47 sn102_47 11.551961
Rsp101_48 sp101_48 sp102_48 11.551961
Rsn101_48 sn101_48 sn102_48 11.551961
Rsp101_49 sp101_49 sp102_49 11.551961
Rsn101_49 sn101_49 sn102_49 11.551961
Rsp101_50 sp101_50 sp102_50 11.551961
Rsn101_50 sn101_50 sn102_50 11.551961
Rsp101_51 sp101_51 sp102_51 11.551961
Rsn101_51 sn101_51 sn102_51 11.551961
Rsp101_52 sp101_52 sp102_52 11.551961
Rsn101_52 sn101_52 sn102_52 11.551961
Rsp101_53 sp101_53 sp102_53 11.551961
Rsn101_53 sn101_53 sn102_53 11.551961
Rsp101_54 sp101_54 sp102_54 11.551961
Rsn101_54 sn101_54 sn102_54 11.551961
Rsp101_55 sp101_55 sp102_55 11.551961
Rsn101_55 sn101_55 sn102_55 11.551961
Rsp101_56 sp101_56 sp102_56 11.551961
Rsn101_56 sn101_56 sn102_56 11.551961
Rsp101_57 sp101_57 sp102_57 11.551961
Rsn101_57 sn101_57 sn102_57 11.551961
Rsp101_58 sp101_58 sp102_58 11.551961
Rsn101_58 sn101_58 sn102_58 11.551961
Rsp101_59 sp101_59 sp102_59 11.551961
Rsn101_59 sn101_59 sn102_59 11.551961
Rsp101_60 sp101_60 sp102_60 11.551961
Rsn101_60 sn101_60 sn102_60 11.551961
Rsp101_61 sp101_61 sp102_61 11.551961
Rsn101_61 sn101_61 sn102_61 11.551961
Rsp101_62 sp101_62 sp102_62 11.551961
Rsn101_62 sn101_62 sn102_62 11.551961
Rsp101_63 sp101_63 sp102_63 11.551961
Rsn101_63 sn101_63 sn102_63 11.551961
Rsp101_64 sp101_64 sp102_64 11.551961
Rsn101_64 sn101_64 sn102_64 11.551961
Rsp101_65 sp101_65 sp102_65 11.551961
Rsn101_65 sn101_65 sn102_65 11.551961
Rsp101_66 sp101_66 sp102_66 11.551961
Rsn101_66 sn101_66 sn102_66 11.551961
Rsp101_67 sp101_67 sp102_67 11.551961
Rsn101_67 sn101_67 sn102_67 11.551961
Rsp101_68 sp101_68 sp102_68 11.551961
Rsn101_68 sn101_68 sn102_68 11.551961
Rsp101_69 sp101_69 sp102_69 11.551961
Rsn101_69 sn101_69 sn102_69 11.551961
Rsp101_70 sp101_70 sp102_70 11.551961
Rsn101_70 sn101_70 sn102_70 11.551961
Rsp101_71 sp101_71 sp102_71 11.551961
Rsn101_71 sn101_71 sn102_71 11.551961
Rsp101_72 sp101_72 sp102_72 11.551961
Rsn101_72 sn101_72 sn102_72 11.551961
Rsp101_73 sp101_73 sp102_73 11.551961
Rsn101_73 sn101_73 sn102_73 11.551961
Rsp101_74 sp101_74 sp102_74 11.551961
Rsn101_74 sn101_74 sn102_74 11.551961
Rsp101_75 sp101_75 sp102_75 11.551961
Rsn101_75 sn101_75 sn102_75 11.551961
Rsp101_76 sp101_76 sp102_76 11.551961
Rsn101_76 sn101_76 sn102_76 11.551961
Rsp101_77 sp101_77 sp102_77 11.551961
Rsn101_77 sn101_77 sn102_77 11.551961
Rsp101_78 sp101_78 sp102_78 11.551961
Rsn101_78 sn101_78 sn102_78 11.551961
Rsp101_79 sp101_79 sp102_79 11.551961
Rsn101_79 sn101_79 sn102_79 11.551961
Rsp101_80 sp101_80 sp102_80 11.551961
Rsn101_80 sn101_80 sn102_80 11.551961
Rsp101_81 sp101_81 sp102_81 11.551961
Rsn101_81 sn101_81 sn102_81 11.551961
Rsp101_82 sp101_82 sp102_82 11.551961
Rsn101_82 sn101_82 sn102_82 11.551961
Rsp101_83 sp101_83 sp102_83 11.551961
Rsn101_83 sn101_83 sn102_83 11.551961
Rsp101_84 sp101_84 sp102_84 11.551961
Rsn101_84 sn101_84 sn102_84 11.551961
Rsp102_1 sp102_1 sp103_1 11.551961
Rsn102_1 sn102_1 sn103_1 11.551961
Rsp102_2 sp102_2 sp103_2 11.551961
Rsn102_2 sn102_2 sn103_2 11.551961
Rsp102_3 sp102_3 sp103_3 11.551961
Rsn102_3 sn102_3 sn103_3 11.551961
Rsp102_4 sp102_4 sp103_4 11.551961
Rsn102_4 sn102_4 sn103_4 11.551961
Rsp102_5 sp102_5 sp103_5 11.551961
Rsn102_5 sn102_5 sn103_5 11.551961
Rsp102_6 sp102_6 sp103_6 11.551961
Rsn102_6 sn102_6 sn103_6 11.551961
Rsp102_7 sp102_7 sp103_7 11.551961
Rsn102_7 sn102_7 sn103_7 11.551961
Rsp102_8 sp102_8 sp103_8 11.551961
Rsn102_8 sn102_8 sn103_8 11.551961
Rsp102_9 sp102_9 sp103_9 11.551961
Rsn102_9 sn102_9 sn103_9 11.551961
Rsp102_10 sp102_10 sp103_10 11.551961
Rsn102_10 sn102_10 sn103_10 11.551961
Rsp102_11 sp102_11 sp103_11 11.551961
Rsn102_11 sn102_11 sn103_11 11.551961
Rsp102_12 sp102_12 sp103_12 11.551961
Rsn102_12 sn102_12 sn103_12 11.551961
Rsp102_13 sp102_13 sp103_13 11.551961
Rsn102_13 sn102_13 sn103_13 11.551961
Rsp102_14 sp102_14 sp103_14 11.551961
Rsn102_14 sn102_14 sn103_14 11.551961
Rsp102_15 sp102_15 sp103_15 11.551961
Rsn102_15 sn102_15 sn103_15 11.551961
Rsp102_16 sp102_16 sp103_16 11.551961
Rsn102_16 sn102_16 sn103_16 11.551961
Rsp102_17 sp102_17 sp103_17 11.551961
Rsn102_17 sn102_17 sn103_17 11.551961
Rsp102_18 sp102_18 sp103_18 11.551961
Rsn102_18 sn102_18 sn103_18 11.551961
Rsp102_19 sp102_19 sp103_19 11.551961
Rsn102_19 sn102_19 sn103_19 11.551961
Rsp102_20 sp102_20 sp103_20 11.551961
Rsn102_20 sn102_20 sn103_20 11.551961
Rsp102_21 sp102_21 sp103_21 11.551961
Rsn102_21 sn102_21 sn103_21 11.551961
Rsp102_22 sp102_22 sp103_22 11.551961
Rsn102_22 sn102_22 sn103_22 11.551961
Rsp102_23 sp102_23 sp103_23 11.551961
Rsn102_23 sn102_23 sn103_23 11.551961
Rsp102_24 sp102_24 sp103_24 11.551961
Rsn102_24 sn102_24 sn103_24 11.551961
Rsp102_25 sp102_25 sp103_25 11.551961
Rsn102_25 sn102_25 sn103_25 11.551961
Rsp102_26 sp102_26 sp103_26 11.551961
Rsn102_26 sn102_26 sn103_26 11.551961
Rsp102_27 sp102_27 sp103_27 11.551961
Rsn102_27 sn102_27 sn103_27 11.551961
Rsp102_28 sp102_28 sp103_28 11.551961
Rsn102_28 sn102_28 sn103_28 11.551961
Rsp102_29 sp102_29 sp103_29 11.551961
Rsn102_29 sn102_29 sn103_29 11.551961
Rsp102_30 sp102_30 sp103_30 11.551961
Rsn102_30 sn102_30 sn103_30 11.551961
Rsp102_31 sp102_31 sp103_31 11.551961
Rsn102_31 sn102_31 sn103_31 11.551961
Rsp102_32 sp102_32 sp103_32 11.551961
Rsn102_32 sn102_32 sn103_32 11.551961
Rsp102_33 sp102_33 sp103_33 11.551961
Rsn102_33 sn102_33 sn103_33 11.551961
Rsp102_34 sp102_34 sp103_34 11.551961
Rsn102_34 sn102_34 sn103_34 11.551961
Rsp102_35 sp102_35 sp103_35 11.551961
Rsn102_35 sn102_35 sn103_35 11.551961
Rsp102_36 sp102_36 sp103_36 11.551961
Rsn102_36 sn102_36 sn103_36 11.551961
Rsp102_37 sp102_37 sp103_37 11.551961
Rsn102_37 sn102_37 sn103_37 11.551961
Rsp102_38 sp102_38 sp103_38 11.551961
Rsn102_38 sn102_38 sn103_38 11.551961
Rsp102_39 sp102_39 sp103_39 11.551961
Rsn102_39 sn102_39 sn103_39 11.551961
Rsp102_40 sp102_40 sp103_40 11.551961
Rsn102_40 sn102_40 sn103_40 11.551961
Rsp102_41 sp102_41 sp103_41 11.551961
Rsn102_41 sn102_41 sn103_41 11.551961
Rsp102_42 sp102_42 sp103_42 11.551961
Rsn102_42 sn102_42 sn103_42 11.551961
Rsp102_43 sp102_43 sp103_43 11.551961
Rsn102_43 sn102_43 sn103_43 11.551961
Rsp102_44 sp102_44 sp103_44 11.551961
Rsn102_44 sn102_44 sn103_44 11.551961
Rsp102_45 sp102_45 sp103_45 11.551961
Rsn102_45 sn102_45 sn103_45 11.551961
Rsp102_46 sp102_46 sp103_46 11.551961
Rsn102_46 sn102_46 sn103_46 11.551961
Rsp102_47 sp102_47 sp103_47 11.551961
Rsn102_47 sn102_47 sn103_47 11.551961
Rsp102_48 sp102_48 sp103_48 11.551961
Rsn102_48 sn102_48 sn103_48 11.551961
Rsp102_49 sp102_49 sp103_49 11.551961
Rsn102_49 sn102_49 sn103_49 11.551961
Rsp102_50 sp102_50 sp103_50 11.551961
Rsn102_50 sn102_50 sn103_50 11.551961
Rsp102_51 sp102_51 sp103_51 11.551961
Rsn102_51 sn102_51 sn103_51 11.551961
Rsp102_52 sp102_52 sp103_52 11.551961
Rsn102_52 sn102_52 sn103_52 11.551961
Rsp102_53 sp102_53 sp103_53 11.551961
Rsn102_53 sn102_53 sn103_53 11.551961
Rsp102_54 sp102_54 sp103_54 11.551961
Rsn102_54 sn102_54 sn103_54 11.551961
Rsp102_55 sp102_55 sp103_55 11.551961
Rsn102_55 sn102_55 sn103_55 11.551961
Rsp102_56 sp102_56 sp103_56 11.551961
Rsn102_56 sn102_56 sn103_56 11.551961
Rsp102_57 sp102_57 sp103_57 11.551961
Rsn102_57 sn102_57 sn103_57 11.551961
Rsp102_58 sp102_58 sp103_58 11.551961
Rsn102_58 sn102_58 sn103_58 11.551961
Rsp102_59 sp102_59 sp103_59 11.551961
Rsn102_59 sn102_59 sn103_59 11.551961
Rsp102_60 sp102_60 sp103_60 11.551961
Rsn102_60 sn102_60 sn103_60 11.551961
Rsp102_61 sp102_61 sp103_61 11.551961
Rsn102_61 sn102_61 sn103_61 11.551961
Rsp102_62 sp102_62 sp103_62 11.551961
Rsn102_62 sn102_62 sn103_62 11.551961
Rsp102_63 sp102_63 sp103_63 11.551961
Rsn102_63 sn102_63 sn103_63 11.551961
Rsp102_64 sp102_64 sp103_64 11.551961
Rsn102_64 sn102_64 sn103_64 11.551961
Rsp102_65 sp102_65 sp103_65 11.551961
Rsn102_65 sn102_65 sn103_65 11.551961
Rsp102_66 sp102_66 sp103_66 11.551961
Rsn102_66 sn102_66 sn103_66 11.551961
Rsp102_67 sp102_67 sp103_67 11.551961
Rsn102_67 sn102_67 sn103_67 11.551961
Rsp102_68 sp102_68 sp103_68 11.551961
Rsn102_68 sn102_68 sn103_68 11.551961
Rsp102_69 sp102_69 sp103_69 11.551961
Rsn102_69 sn102_69 sn103_69 11.551961
Rsp102_70 sp102_70 sp103_70 11.551961
Rsn102_70 sn102_70 sn103_70 11.551961
Rsp102_71 sp102_71 sp103_71 11.551961
Rsn102_71 sn102_71 sn103_71 11.551961
Rsp102_72 sp102_72 sp103_72 11.551961
Rsn102_72 sn102_72 sn103_72 11.551961
Rsp102_73 sp102_73 sp103_73 11.551961
Rsn102_73 sn102_73 sn103_73 11.551961
Rsp102_74 sp102_74 sp103_74 11.551961
Rsn102_74 sn102_74 sn103_74 11.551961
Rsp102_75 sp102_75 sp103_75 11.551961
Rsn102_75 sn102_75 sn103_75 11.551961
Rsp102_76 sp102_76 sp103_76 11.551961
Rsn102_76 sn102_76 sn103_76 11.551961
Rsp102_77 sp102_77 sp103_77 11.551961
Rsn102_77 sn102_77 sn103_77 11.551961
Rsp102_78 sp102_78 sp103_78 11.551961
Rsn102_78 sn102_78 sn103_78 11.551961
Rsp102_79 sp102_79 sp103_79 11.551961
Rsn102_79 sn102_79 sn103_79 11.551961
Rsp102_80 sp102_80 sp103_80 11.551961
Rsn102_80 sn102_80 sn103_80 11.551961
Rsp102_81 sp102_81 sp103_81 11.551961
Rsn102_81 sn102_81 sn103_81 11.551961
Rsp102_82 sp102_82 sp103_82 11.551961
Rsn102_82 sn102_82 sn103_82 11.551961
Rsp102_83 sp102_83 sp103_83 11.551961
Rsn102_83 sn102_83 sn103_83 11.551961
Rsp102_84 sp102_84 sp103_84 11.551961
Rsn102_84 sn102_84 sn103_84 11.551961
Rsp103_1 sp103_1 sp104_1 11.551961
Rsn103_1 sn103_1 sn104_1 11.551961
Rsp103_2 sp103_2 sp104_2 11.551961
Rsn103_2 sn103_2 sn104_2 11.551961
Rsp103_3 sp103_3 sp104_3 11.551961
Rsn103_3 sn103_3 sn104_3 11.551961
Rsp103_4 sp103_4 sp104_4 11.551961
Rsn103_4 sn103_4 sn104_4 11.551961
Rsp103_5 sp103_5 sp104_5 11.551961
Rsn103_5 sn103_5 sn104_5 11.551961
Rsp103_6 sp103_6 sp104_6 11.551961
Rsn103_6 sn103_6 sn104_6 11.551961
Rsp103_7 sp103_7 sp104_7 11.551961
Rsn103_7 sn103_7 sn104_7 11.551961
Rsp103_8 sp103_8 sp104_8 11.551961
Rsn103_8 sn103_8 sn104_8 11.551961
Rsp103_9 sp103_9 sp104_9 11.551961
Rsn103_9 sn103_9 sn104_9 11.551961
Rsp103_10 sp103_10 sp104_10 11.551961
Rsn103_10 sn103_10 sn104_10 11.551961
Rsp103_11 sp103_11 sp104_11 11.551961
Rsn103_11 sn103_11 sn104_11 11.551961
Rsp103_12 sp103_12 sp104_12 11.551961
Rsn103_12 sn103_12 sn104_12 11.551961
Rsp103_13 sp103_13 sp104_13 11.551961
Rsn103_13 sn103_13 sn104_13 11.551961
Rsp103_14 sp103_14 sp104_14 11.551961
Rsn103_14 sn103_14 sn104_14 11.551961
Rsp103_15 sp103_15 sp104_15 11.551961
Rsn103_15 sn103_15 sn104_15 11.551961
Rsp103_16 sp103_16 sp104_16 11.551961
Rsn103_16 sn103_16 sn104_16 11.551961
Rsp103_17 sp103_17 sp104_17 11.551961
Rsn103_17 sn103_17 sn104_17 11.551961
Rsp103_18 sp103_18 sp104_18 11.551961
Rsn103_18 sn103_18 sn104_18 11.551961
Rsp103_19 sp103_19 sp104_19 11.551961
Rsn103_19 sn103_19 sn104_19 11.551961
Rsp103_20 sp103_20 sp104_20 11.551961
Rsn103_20 sn103_20 sn104_20 11.551961
Rsp103_21 sp103_21 sp104_21 11.551961
Rsn103_21 sn103_21 sn104_21 11.551961
Rsp103_22 sp103_22 sp104_22 11.551961
Rsn103_22 sn103_22 sn104_22 11.551961
Rsp103_23 sp103_23 sp104_23 11.551961
Rsn103_23 sn103_23 sn104_23 11.551961
Rsp103_24 sp103_24 sp104_24 11.551961
Rsn103_24 sn103_24 sn104_24 11.551961
Rsp103_25 sp103_25 sp104_25 11.551961
Rsn103_25 sn103_25 sn104_25 11.551961
Rsp103_26 sp103_26 sp104_26 11.551961
Rsn103_26 sn103_26 sn104_26 11.551961
Rsp103_27 sp103_27 sp104_27 11.551961
Rsn103_27 sn103_27 sn104_27 11.551961
Rsp103_28 sp103_28 sp104_28 11.551961
Rsn103_28 sn103_28 sn104_28 11.551961
Rsp103_29 sp103_29 sp104_29 11.551961
Rsn103_29 sn103_29 sn104_29 11.551961
Rsp103_30 sp103_30 sp104_30 11.551961
Rsn103_30 sn103_30 sn104_30 11.551961
Rsp103_31 sp103_31 sp104_31 11.551961
Rsn103_31 sn103_31 sn104_31 11.551961
Rsp103_32 sp103_32 sp104_32 11.551961
Rsn103_32 sn103_32 sn104_32 11.551961
Rsp103_33 sp103_33 sp104_33 11.551961
Rsn103_33 sn103_33 sn104_33 11.551961
Rsp103_34 sp103_34 sp104_34 11.551961
Rsn103_34 sn103_34 sn104_34 11.551961
Rsp103_35 sp103_35 sp104_35 11.551961
Rsn103_35 sn103_35 sn104_35 11.551961
Rsp103_36 sp103_36 sp104_36 11.551961
Rsn103_36 sn103_36 sn104_36 11.551961
Rsp103_37 sp103_37 sp104_37 11.551961
Rsn103_37 sn103_37 sn104_37 11.551961
Rsp103_38 sp103_38 sp104_38 11.551961
Rsn103_38 sn103_38 sn104_38 11.551961
Rsp103_39 sp103_39 sp104_39 11.551961
Rsn103_39 sn103_39 sn104_39 11.551961
Rsp103_40 sp103_40 sp104_40 11.551961
Rsn103_40 sn103_40 sn104_40 11.551961
Rsp103_41 sp103_41 sp104_41 11.551961
Rsn103_41 sn103_41 sn104_41 11.551961
Rsp103_42 sp103_42 sp104_42 11.551961
Rsn103_42 sn103_42 sn104_42 11.551961
Rsp103_43 sp103_43 sp104_43 11.551961
Rsn103_43 sn103_43 sn104_43 11.551961
Rsp103_44 sp103_44 sp104_44 11.551961
Rsn103_44 sn103_44 sn104_44 11.551961
Rsp103_45 sp103_45 sp104_45 11.551961
Rsn103_45 sn103_45 sn104_45 11.551961
Rsp103_46 sp103_46 sp104_46 11.551961
Rsn103_46 sn103_46 sn104_46 11.551961
Rsp103_47 sp103_47 sp104_47 11.551961
Rsn103_47 sn103_47 sn104_47 11.551961
Rsp103_48 sp103_48 sp104_48 11.551961
Rsn103_48 sn103_48 sn104_48 11.551961
Rsp103_49 sp103_49 sp104_49 11.551961
Rsn103_49 sn103_49 sn104_49 11.551961
Rsp103_50 sp103_50 sp104_50 11.551961
Rsn103_50 sn103_50 sn104_50 11.551961
Rsp103_51 sp103_51 sp104_51 11.551961
Rsn103_51 sn103_51 sn104_51 11.551961
Rsp103_52 sp103_52 sp104_52 11.551961
Rsn103_52 sn103_52 sn104_52 11.551961
Rsp103_53 sp103_53 sp104_53 11.551961
Rsn103_53 sn103_53 sn104_53 11.551961
Rsp103_54 sp103_54 sp104_54 11.551961
Rsn103_54 sn103_54 sn104_54 11.551961
Rsp103_55 sp103_55 sp104_55 11.551961
Rsn103_55 sn103_55 sn104_55 11.551961
Rsp103_56 sp103_56 sp104_56 11.551961
Rsn103_56 sn103_56 sn104_56 11.551961
Rsp103_57 sp103_57 sp104_57 11.551961
Rsn103_57 sn103_57 sn104_57 11.551961
Rsp103_58 sp103_58 sp104_58 11.551961
Rsn103_58 sn103_58 sn104_58 11.551961
Rsp103_59 sp103_59 sp104_59 11.551961
Rsn103_59 sn103_59 sn104_59 11.551961
Rsp103_60 sp103_60 sp104_60 11.551961
Rsn103_60 sn103_60 sn104_60 11.551961
Rsp103_61 sp103_61 sp104_61 11.551961
Rsn103_61 sn103_61 sn104_61 11.551961
Rsp103_62 sp103_62 sp104_62 11.551961
Rsn103_62 sn103_62 sn104_62 11.551961
Rsp103_63 sp103_63 sp104_63 11.551961
Rsn103_63 sn103_63 sn104_63 11.551961
Rsp103_64 sp103_64 sp104_64 11.551961
Rsn103_64 sn103_64 sn104_64 11.551961
Rsp103_65 sp103_65 sp104_65 11.551961
Rsn103_65 sn103_65 sn104_65 11.551961
Rsp103_66 sp103_66 sp104_66 11.551961
Rsn103_66 sn103_66 sn104_66 11.551961
Rsp103_67 sp103_67 sp104_67 11.551961
Rsn103_67 sn103_67 sn104_67 11.551961
Rsp103_68 sp103_68 sp104_68 11.551961
Rsn103_68 sn103_68 sn104_68 11.551961
Rsp103_69 sp103_69 sp104_69 11.551961
Rsn103_69 sn103_69 sn104_69 11.551961
Rsp103_70 sp103_70 sp104_70 11.551961
Rsn103_70 sn103_70 sn104_70 11.551961
Rsp103_71 sp103_71 sp104_71 11.551961
Rsn103_71 sn103_71 sn104_71 11.551961
Rsp103_72 sp103_72 sp104_72 11.551961
Rsn103_72 sn103_72 sn104_72 11.551961
Rsp103_73 sp103_73 sp104_73 11.551961
Rsn103_73 sn103_73 sn104_73 11.551961
Rsp103_74 sp103_74 sp104_74 11.551961
Rsn103_74 sn103_74 sn104_74 11.551961
Rsp103_75 sp103_75 sp104_75 11.551961
Rsn103_75 sn103_75 sn104_75 11.551961
Rsp103_76 sp103_76 sp104_76 11.551961
Rsn103_76 sn103_76 sn104_76 11.551961
Rsp103_77 sp103_77 sp104_77 11.551961
Rsn103_77 sn103_77 sn104_77 11.551961
Rsp103_78 sp103_78 sp104_78 11.551961
Rsn103_78 sn103_78 sn104_78 11.551961
Rsp103_79 sp103_79 sp104_79 11.551961
Rsn103_79 sn103_79 sn104_79 11.551961
Rsp103_80 sp103_80 sp104_80 11.551961
Rsn103_80 sn103_80 sn104_80 11.551961
Rsp103_81 sp103_81 sp104_81 11.551961
Rsn103_81 sn103_81 sn104_81 11.551961
Rsp103_82 sp103_82 sp104_82 11.551961
Rsn103_82 sn103_82 sn104_82 11.551961
Rsp103_83 sp103_83 sp104_83 11.551961
Rsn103_83 sn103_83 sn104_83 11.551961
Rsp103_84 sp103_84 sp104_84 11.551961
Rsn103_84 sn103_84 sn104_84 11.551961
Rsp104_1 sp104_1 sp105_1 11.551961
Rsn104_1 sn104_1 sn105_1 11.551961
Rsp104_2 sp104_2 sp105_2 11.551961
Rsn104_2 sn104_2 sn105_2 11.551961
Rsp104_3 sp104_3 sp105_3 11.551961
Rsn104_3 sn104_3 sn105_3 11.551961
Rsp104_4 sp104_4 sp105_4 11.551961
Rsn104_4 sn104_4 sn105_4 11.551961
Rsp104_5 sp104_5 sp105_5 11.551961
Rsn104_5 sn104_5 sn105_5 11.551961
Rsp104_6 sp104_6 sp105_6 11.551961
Rsn104_6 sn104_6 sn105_6 11.551961
Rsp104_7 sp104_7 sp105_7 11.551961
Rsn104_7 sn104_7 sn105_7 11.551961
Rsp104_8 sp104_8 sp105_8 11.551961
Rsn104_8 sn104_8 sn105_8 11.551961
Rsp104_9 sp104_9 sp105_9 11.551961
Rsn104_9 sn104_9 sn105_9 11.551961
Rsp104_10 sp104_10 sp105_10 11.551961
Rsn104_10 sn104_10 sn105_10 11.551961
Rsp104_11 sp104_11 sp105_11 11.551961
Rsn104_11 sn104_11 sn105_11 11.551961
Rsp104_12 sp104_12 sp105_12 11.551961
Rsn104_12 sn104_12 sn105_12 11.551961
Rsp104_13 sp104_13 sp105_13 11.551961
Rsn104_13 sn104_13 sn105_13 11.551961
Rsp104_14 sp104_14 sp105_14 11.551961
Rsn104_14 sn104_14 sn105_14 11.551961
Rsp104_15 sp104_15 sp105_15 11.551961
Rsn104_15 sn104_15 sn105_15 11.551961
Rsp104_16 sp104_16 sp105_16 11.551961
Rsn104_16 sn104_16 sn105_16 11.551961
Rsp104_17 sp104_17 sp105_17 11.551961
Rsn104_17 sn104_17 sn105_17 11.551961
Rsp104_18 sp104_18 sp105_18 11.551961
Rsn104_18 sn104_18 sn105_18 11.551961
Rsp104_19 sp104_19 sp105_19 11.551961
Rsn104_19 sn104_19 sn105_19 11.551961
Rsp104_20 sp104_20 sp105_20 11.551961
Rsn104_20 sn104_20 sn105_20 11.551961
Rsp104_21 sp104_21 sp105_21 11.551961
Rsn104_21 sn104_21 sn105_21 11.551961
Rsp104_22 sp104_22 sp105_22 11.551961
Rsn104_22 sn104_22 sn105_22 11.551961
Rsp104_23 sp104_23 sp105_23 11.551961
Rsn104_23 sn104_23 sn105_23 11.551961
Rsp104_24 sp104_24 sp105_24 11.551961
Rsn104_24 sn104_24 sn105_24 11.551961
Rsp104_25 sp104_25 sp105_25 11.551961
Rsn104_25 sn104_25 sn105_25 11.551961
Rsp104_26 sp104_26 sp105_26 11.551961
Rsn104_26 sn104_26 sn105_26 11.551961
Rsp104_27 sp104_27 sp105_27 11.551961
Rsn104_27 sn104_27 sn105_27 11.551961
Rsp104_28 sp104_28 sp105_28 11.551961
Rsn104_28 sn104_28 sn105_28 11.551961
Rsp104_29 sp104_29 sp105_29 11.551961
Rsn104_29 sn104_29 sn105_29 11.551961
Rsp104_30 sp104_30 sp105_30 11.551961
Rsn104_30 sn104_30 sn105_30 11.551961
Rsp104_31 sp104_31 sp105_31 11.551961
Rsn104_31 sn104_31 sn105_31 11.551961
Rsp104_32 sp104_32 sp105_32 11.551961
Rsn104_32 sn104_32 sn105_32 11.551961
Rsp104_33 sp104_33 sp105_33 11.551961
Rsn104_33 sn104_33 sn105_33 11.551961
Rsp104_34 sp104_34 sp105_34 11.551961
Rsn104_34 sn104_34 sn105_34 11.551961
Rsp104_35 sp104_35 sp105_35 11.551961
Rsn104_35 sn104_35 sn105_35 11.551961
Rsp104_36 sp104_36 sp105_36 11.551961
Rsn104_36 sn104_36 sn105_36 11.551961
Rsp104_37 sp104_37 sp105_37 11.551961
Rsn104_37 sn104_37 sn105_37 11.551961
Rsp104_38 sp104_38 sp105_38 11.551961
Rsn104_38 sn104_38 sn105_38 11.551961
Rsp104_39 sp104_39 sp105_39 11.551961
Rsn104_39 sn104_39 sn105_39 11.551961
Rsp104_40 sp104_40 sp105_40 11.551961
Rsn104_40 sn104_40 sn105_40 11.551961
Rsp104_41 sp104_41 sp105_41 11.551961
Rsn104_41 sn104_41 sn105_41 11.551961
Rsp104_42 sp104_42 sp105_42 11.551961
Rsn104_42 sn104_42 sn105_42 11.551961
Rsp104_43 sp104_43 sp105_43 11.551961
Rsn104_43 sn104_43 sn105_43 11.551961
Rsp104_44 sp104_44 sp105_44 11.551961
Rsn104_44 sn104_44 sn105_44 11.551961
Rsp104_45 sp104_45 sp105_45 11.551961
Rsn104_45 sn104_45 sn105_45 11.551961
Rsp104_46 sp104_46 sp105_46 11.551961
Rsn104_46 sn104_46 sn105_46 11.551961
Rsp104_47 sp104_47 sp105_47 11.551961
Rsn104_47 sn104_47 sn105_47 11.551961
Rsp104_48 sp104_48 sp105_48 11.551961
Rsn104_48 sn104_48 sn105_48 11.551961
Rsp104_49 sp104_49 sp105_49 11.551961
Rsn104_49 sn104_49 sn105_49 11.551961
Rsp104_50 sp104_50 sp105_50 11.551961
Rsn104_50 sn104_50 sn105_50 11.551961
Rsp104_51 sp104_51 sp105_51 11.551961
Rsn104_51 sn104_51 sn105_51 11.551961
Rsp104_52 sp104_52 sp105_52 11.551961
Rsn104_52 sn104_52 sn105_52 11.551961
Rsp104_53 sp104_53 sp105_53 11.551961
Rsn104_53 sn104_53 sn105_53 11.551961
Rsp104_54 sp104_54 sp105_54 11.551961
Rsn104_54 sn104_54 sn105_54 11.551961
Rsp104_55 sp104_55 sp105_55 11.551961
Rsn104_55 sn104_55 sn105_55 11.551961
Rsp104_56 sp104_56 sp105_56 11.551961
Rsn104_56 sn104_56 sn105_56 11.551961
Rsp104_57 sp104_57 sp105_57 11.551961
Rsn104_57 sn104_57 sn105_57 11.551961
Rsp104_58 sp104_58 sp105_58 11.551961
Rsn104_58 sn104_58 sn105_58 11.551961
Rsp104_59 sp104_59 sp105_59 11.551961
Rsn104_59 sn104_59 sn105_59 11.551961
Rsp104_60 sp104_60 sp105_60 11.551961
Rsn104_60 sn104_60 sn105_60 11.551961
Rsp104_61 sp104_61 sp105_61 11.551961
Rsn104_61 sn104_61 sn105_61 11.551961
Rsp104_62 sp104_62 sp105_62 11.551961
Rsn104_62 sn104_62 sn105_62 11.551961
Rsp104_63 sp104_63 sp105_63 11.551961
Rsn104_63 sn104_63 sn105_63 11.551961
Rsp104_64 sp104_64 sp105_64 11.551961
Rsn104_64 sn104_64 sn105_64 11.551961
Rsp104_65 sp104_65 sp105_65 11.551961
Rsn104_65 sn104_65 sn105_65 11.551961
Rsp104_66 sp104_66 sp105_66 11.551961
Rsn104_66 sn104_66 sn105_66 11.551961
Rsp104_67 sp104_67 sp105_67 11.551961
Rsn104_67 sn104_67 sn105_67 11.551961
Rsp104_68 sp104_68 sp105_68 11.551961
Rsn104_68 sn104_68 sn105_68 11.551961
Rsp104_69 sp104_69 sp105_69 11.551961
Rsn104_69 sn104_69 sn105_69 11.551961
Rsp104_70 sp104_70 sp105_70 11.551961
Rsn104_70 sn104_70 sn105_70 11.551961
Rsp104_71 sp104_71 sp105_71 11.551961
Rsn104_71 sn104_71 sn105_71 11.551961
Rsp104_72 sp104_72 sp105_72 11.551961
Rsn104_72 sn104_72 sn105_72 11.551961
Rsp104_73 sp104_73 sp105_73 11.551961
Rsn104_73 sn104_73 sn105_73 11.551961
Rsp104_74 sp104_74 sp105_74 11.551961
Rsn104_74 sn104_74 sn105_74 11.551961
Rsp104_75 sp104_75 sp105_75 11.551961
Rsn104_75 sn104_75 sn105_75 11.551961
Rsp104_76 sp104_76 sp105_76 11.551961
Rsn104_76 sn104_76 sn105_76 11.551961
Rsp104_77 sp104_77 sp105_77 11.551961
Rsn104_77 sn104_77 sn105_77 11.551961
Rsp104_78 sp104_78 sp105_78 11.551961
Rsn104_78 sn104_78 sn105_78 11.551961
Rsp104_79 sp104_79 sp105_79 11.551961
Rsn104_79 sn104_79 sn105_79 11.551961
Rsp104_80 sp104_80 sp105_80 11.551961
Rsn104_80 sn104_80 sn105_80 11.551961
Rsp104_81 sp104_81 sp105_81 11.551961
Rsn104_81 sn104_81 sn105_81 11.551961
Rsp104_82 sp104_82 sp105_82 11.551961
Rsn104_82 sn104_82 sn105_82 11.551961
Rsp104_83 sp104_83 sp105_83 11.551961
Rsn104_83 sn104_83 sn105_83 11.551961
Rsp104_84 sp104_84 sp105_84 11.551961
Rsn104_84 sn104_84 sn105_84 11.551961
Rsp105_1 sp105_1 sp106_1 11.551961
Rsn105_1 sn105_1 sn106_1 11.551961
Rsp105_2 sp105_2 sp106_2 11.551961
Rsn105_2 sn105_2 sn106_2 11.551961
Rsp105_3 sp105_3 sp106_3 11.551961
Rsn105_3 sn105_3 sn106_3 11.551961
Rsp105_4 sp105_4 sp106_4 11.551961
Rsn105_4 sn105_4 sn106_4 11.551961
Rsp105_5 sp105_5 sp106_5 11.551961
Rsn105_5 sn105_5 sn106_5 11.551961
Rsp105_6 sp105_6 sp106_6 11.551961
Rsn105_6 sn105_6 sn106_6 11.551961
Rsp105_7 sp105_7 sp106_7 11.551961
Rsn105_7 sn105_7 sn106_7 11.551961
Rsp105_8 sp105_8 sp106_8 11.551961
Rsn105_8 sn105_8 sn106_8 11.551961
Rsp105_9 sp105_9 sp106_9 11.551961
Rsn105_9 sn105_9 sn106_9 11.551961
Rsp105_10 sp105_10 sp106_10 11.551961
Rsn105_10 sn105_10 sn106_10 11.551961
Rsp105_11 sp105_11 sp106_11 11.551961
Rsn105_11 sn105_11 sn106_11 11.551961
Rsp105_12 sp105_12 sp106_12 11.551961
Rsn105_12 sn105_12 sn106_12 11.551961
Rsp105_13 sp105_13 sp106_13 11.551961
Rsn105_13 sn105_13 sn106_13 11.551961
Rsp105_14 sp105_14 sp106_14 11.551961
Rsn105_14 sn105_14 sn106_14 11.551961
Rsp105_15 sp105_15 sp106_15 11.551961
Rsn105_15 sn105_15 sn106_15 11.551961
Rsp105_16 sp105_16 sp106_16 11.551961
Rsn105_16 sn105_16 sn106_16 11.551961
Rsp105_17 sp105_17 sp106_17 11.551961
Rsn105_17 sn105_17 sn106_17 11.551961
Rsp105_18 sp105_18 sp106_18 11.551961
Rsn105_18 sn105_18 sn106_18 11.551961
Rsp105_19 sp105_19 sp106_19 11.551961
Rsn105_19 sn105_19 sn106_19 11.551961
Rsp105_20 sp105_20 sp106_20 11.551961
Rsn105_20 sn105_20 sn106_20 11.551961
Rsp105_21 sp105_21 sp106_21 11.551961
Rsn105_21 sn105_21 sn106_21 11.551961
Rsp105_22 sp105_22 sp106_22 11.551961
Rsn105_22 sn105_22 sn106_22 11.551961
Rsp105_23 sp105_23 sp106_23 11.551961
Rsn105_23 sn105_23 sn106_23 11.551961
Rsp105_24 sp105_24 sp106_24 11.551961
Rsn105_24 sn105_24 sn106_24 11.551961
Rsp105_25 sp105_25 sp106_25 11.551961
Rsn105_25 sn105_25 sn106_25 11.551961
Rsp105_26 sp105_26 sp106_26 11.551961
Rsn105_26 sn105_26 sn106_26 11.551961
Rsp105_27 sp105_27 sp106_27 11.551961
Rsn105_27 sn105_27 sn106_27 11.551961
Rsp105_28 sp105_28 sp106_28 11.551961
Rsn105_28 sn105_28 sn106_28 11.551961
Rsp105_29 sp105_29 sp106_29 11.551961
Rsn105_29 sn105_29 sn106_29 11.551961
Rsp105_30 sp105_30 sp106_30 11.551961
Rsn105_30 sn105_30 sn106_30 11.551961
Rsp105_31 sp105_31 sp106_31 11.551961
Rsn105_31 sn105_31 sn106_31 11.551961
Rsp105_32 sp105_32 sp106_32 11.551961
Rsn105_32 sn105_32 sn106_32 11.551961
Rsp105_33 sp105_33 sp106_33 11.551961
Rsn105_33 sn105_33 sn106_33 11.551961
Rsp105_34 sp105_34 sp106_34 11.551961
Rsn105_34 sn105_34 sn106_34 11.551961
Rsp105_35 sp105_35 sp106_35 11.551961
Rsn105_35 sn105_35 sn106_35 11.551961
Rsp105_36 sp105_36 sp106_36 11.551961
Rsn105_36 sn105_36 sn106_36 11.551961
Rsp105_37 sp105_37 sp106_37 11.551961
Rsn105_37 sn105_37 sn106_37 11.551961
Rsp105_38 sp105_38 sp106_38 11.551961
Rsn105_38 sn105_38 sn106_38 11.551961
Rsp105_39 sp105_39 sp106_39 11.551961
Rsn105_39 sn105_39 sn106_39 11.551961
Rsp105_40 sp105_40 sp106_40 11.551961
Rsn105_40 sn105_40 sn106_40 11.551961
Rsp105_41 sp105_41 sp106_41 11.551961
Rsn105_41 sn105_41 sn106_41 11.551961
Rsp105_42 sp105_42 sp106_42 11.551961
Rsn105_42 sn105_42 sn106_42 11.551961
Rsp105_43 sp105_43 sp106_43 11.551961
Rsn105_43 sn105_43 sn106_43 11.551961
Rsp105_44 sp105_44 sp106_44 11.551961
Rsn105_44 sn105_44 sn106_44 11.551961
Rsp105_45 sp105_45 sp106_45 11.551961
Rsn105_45 sn105_45 sn106_45 11.551961
Rsp105_46 sp105_46 sp106_46 11.551961
Rsn105_46 sn105_46 sn106_46 11.551961
Rsp105_47 sp105_47 sp106_47 11.551961
Rsn105_47 sn105_47 sn106_47 11.551961
Rsp105_48 sp105_48 sp106_48 11.551961
Rsn105_48 sn105_48 sn106_48 11.551961
Rsp105_49 sp105_49 sp106_49 11.551961
Rsn105_49 sn105_49 sn106_49 11.551961
Rsp105_50 sp105_50 sp106_50 11.551961
Rsn105_50 sn105_50 sn106_50 11.551961
Rsp105_51 sp105_51 sp106_51 11.551961
Rsn105_51 sn105_51 sn106_51 11.551961
Rsp105_52 sp105_52 sp106_52 11.551961
Rsn105_52 sn105_52 sn106_52 11.551961
Rsp105_53 sp105_53 sp106_53 11.551961
Rsn105_53 sn105_53 sn106_53 11.551961
Rsp105_54 sp105_54 sp106_54 11.551961
Rsn105_54 sn105_54 sn106_54 11.551961
Rsp105_55 sp105_55 sp106_55 11.551961
Rsn105_55 sn105_55 sn106_55 11.551961
Rsp105_56 sp105_56 sp106_56 11.551961
Rsn105_56 sn105_56 sn106_56 11.551961
Rsp105_57 sp105_57 sp106_57 11.551961
Rsn105_57 sn105_57 sn106_57 11.551961
Rsp105_58 sp105_58 sp106_58 11.551961
Rsn105_58 sn105_58 sn106_58 11.551961
Rsp105_59 sp105_59 sp106_59 11.551961
Rsn105_59 sn105_59 sn106_59 11.551961
Rsp105_60 sp105_60 sp106_60 11.551961
Rsn105_60 sn105_60 sn106_60 11.551961
Rsp105_61 sp105_61 sp106_61 11.551961
Rsn105_61 sn105_61 sn106_61 11.551961
Rsp105_62 sp105_62 sp106_62 11.551961
Rsn105_62 sn105_62 sn106_62 11.551961
Rsp105_63 sp105_63 sp106_63 11.551961
Rsn105_63 sn105_63 sn106_63 11.551961
Rsp105_64 sp105_64 sp106_64 11.551961
Rsn105_64 sn105_64 sn106_64 11.551961
Rsp105_65 sp105_65 sp106_65 11.551961
Rsn105_65 sn105_65 sn106_65 11.551961
Rsp105_66 sp105_66 sp106_66 11.551961
Rsn105_66 sn105_66 sn106_66 11.551961
Rsp105_67 sp105_67 sp106_67 11.551961
Rsn105_67 sn105_67 sn106_67 11.551961
Rsp105_68 sp105_68 sp106_68 11.551961
Rsn105_68 sn105_68 sn106_68 11.551961
Rsp105_69 sp105_69 sp106_69 11.551961
Rsn105_69 sn105_69 sn106_69 11.551961
Rsp105_70 sp105_70 sp106_70 11.551961
Rsn105_70 sn105_70 sn106_70 11.551961
Rsp105_71 sp105_71 sp106_71 11.551961
Rsn105_71 sn105_71 sn106_71 11.551961
Rsp105_72 sp105_72 sp106_72 11.551961
Rsn105_72 sn105_72 sn106_72 11.551961
Rsp105_73 sp105_73 sp106_73 11.551961
Rsn105_73 sn105_73 sn106_73 11.551961
Rsp105_74 sp105_74 sp106_74 11.551961
Rsn105_74 sn105_74 sn106_74 11.551961
Rsp105_75 sp105_75 sp106_75 11.551961
Rsn105_75 sn105_75 sn106_75 11.551961
Rsp105_76 sp105_76 sp106_76 11.551961
Rsn105_76 sn105_76 sn106_76 11.551961
Rsp105_77 sp105_77 sp106_77 11.551961
Rsn105_77 sn105_77 sn106_77 11.551961
Rsp105_78 sp105_78 sp106_78 11.551961
Rsn105_78 sn105_78 sn106_78 11.551961
Rsp105_79 sp105_79 sp106_79 11.551961
Rsn105_79 sn105_79 sn106_79 11.551961
Rsp105_80 sp105_80 sp106_80 11.551961
Rsn105_80 sn105_80 sn106_80 11.551961
Rsp105_81 sp105_81 sp106_81 11.551961
Rsn105_81 sn105_81 sn106_81 11.551961
Rsp105_82 sp105_82 sp106_82 11.551961
Rsn105_82 sn105_82 sn106_82 11.551961
Rsp105_83 sp105_83 sp106_83 11.551961
Rsn105_83 sn105_83 sn106_83 11.551961
Rsp105_84 sp105_84 sp106_84 11.551961
Rsn105_84 sn105_84 sn106_84 11.551961
Rsp106_1 sp106_1 sp107_1 11.551961
Rsn106_1 sn106_1 sn107_1 11.551961
Rsp106_2 sp106_2 sp107_2 11.551961
Rsn106_2 sn106_2 sn107_2 11.551961
Rsp106_3 sp106_3 sp107_3 11.551961
Rsn106_3 sn106_3 sn107_3 11.551961
Rsp106_4 sp106_4 sp107_4 11.551961
Rsn106_4 sn106_4 sn107_4 11.551961
Rsp106_5 sp106_5 sp107_5 11.551961
Rsn106_5 sn106_5 sn107_5 11.551961
Rsp106_6 sp106_6 sp107_6 11.551961
Rsn106_6 sn106_6 sn107_6 11.551961
Rsp106_7 sp106_7 sp107_7 11.551961
Rsn106_7 sn106_7 sn107_7 11.551961
Rsp106_8 sp106_8 sp107_8 11.551961
Rsn106_8 sn106_8 sn107_8 11.551961
Rsp106_9 sp106_9 sp107_9 11.551961
Rsn106_9 sn106_9 sn107_9 11.551961
Rsp106_10 sp106_10 sp107_10 11.551961
Rsn106_10 sn106_10 sn107_10 11.551961
Rsp106_11 sp106_11 sp107_11 11.551961
Rsn106_11 sn106_11 sn107_11 11.551961
Rsp106_12 sp106_12 sp107_12 11.551961
Rsn106_12 sn106_12 sn107_12 11.551961
Rsp106_13 sp106_13 sp107_13 11.551961
Rsn106_13 sn106_13 sn107_13 11.551961
Rsp106_14 sp106_14 sp107_14 11.551961
Rsn106_14 sn106_14 sn107_14 11.551961
Rsp106_15 sp106_15 sp107_15 11.551961
Rsn106_15 sn106_15 sn107_15 11.551961
Rsp106_16 sp106_16 sp107_16 11.551961
Rsn106_16 sn106_16 sn107_16 11.551961
Rsp106_17 sp106_17 sp107_17 11.551961
Rsn106_17 sn106_17 sn107_17 11.551961
Rsp106_18 sp106_18 sp107_18 11.551961
Rsn106_18 sn106_18 sn107_18 11.551961
Rsp106_19 sp106_19 sp107_19 11.551961
Rsn106_19 sn106_19 sn107_19 11.551961
Rsp106_20 sp106_20 sp107_20 11.551961
Rsn106_20 sn106_20 sn107_20 11.551961
Rsp106_21 sp106_21 sp107_21 11.551961
Rsn106_21 sn106_21 sn107_21 11.551961
Rsp106_22 sp106_22 sp107_22 11.551961
Rsn106_22 sn106_22 sn107_22 11.551961
Rsp106_23 sp106_23 sp107_23 11.551961
Rsn106_23 sn106_23 sn107_23 11.551961
Rsp106_24 sp106_24 sp107_24 11.551961
Rsn106_24 sn106_24 sn107_24 11.551961
Rsp106_25 sp106_25 sp107_25 11.551961
Rsn106_25 sn106_25 sn107_25 11.551961
Rsp106_26 sp106_26 sp107_26 11.551961
Rsn106_26 sn106_26 sn107_26 11.551961
Rsp106_27 sp106_27 sp107_27 11.551961
Rsn106_27 sn106_27 sn107_27 11.551961
Rsp106_28 sp106_28 sp107_28 11.551961
Rsn106_28 sn106_28 sn107_28 11.551961
Rsp106_29 sp106_29 sp107_29 11.551961
Rsn106_29 sn106_29 sn107_29 11.551961
Rsp106_30 sp106_30 sp107_30 11.551961
Rsn106_30 sn106_30 sn107_30 11.551961
Rsp106_31 sp106_31 sp107_31 11.551961
Rsn106_31 sn106_31 sn107_31 11.551961
Rsp106_32 sp106_32 sp107_32 11.551961
Rsn106_32 sn106_32 sn107_32 11.551961
Rsp106_33 sp106_33 sp107_33 11.551961
Rsn106_33 sn106_33 sn107_33 11.551961
Rsp106_34 sp106_34 sp107_34 11.551961
Rsn106_34 sn106_34 sn107_34 11.551961
Rsp106_35 sp106_35 sp107_35 11.551961
Rsn106_35 sn106_35 sn107_35 11.551961
Rsp106_36 sp106_36 sp107_36 11.551961
Rsn106_36 sn106_36 sn107_36 11.551961
Rsp106_37 sp106_37 sp107_37 11.551961
Rsn106_37 sn106_37 sn107_37 11.551961
Rsp106_38 sp106_38 sp107_38 11.551961
Rsn106_38 sn106_38 sn107_38 11.551961
Rsp106_39 sp106_39 sp107_39 11.551961
Rsn106_39 sn106_39 sn107_39 11.551961
Rsp106_40 sp106_40 sp107_40 11.551961
Rsn106_40 sn106_40 sn107_40 11.551961
Rsp106_41 sp106_41 sp107_41 11.551961
Rsn106_41 sn106_41 sn107_41 11.551961
Rsp106_42 sp106_42 sp107_42 11.551961
Rsn106_42 sn106_42 sn107_42 11.551961
Rsp106_43 sp106_43 sp107_43 11.551961
Rsn106_43 sn106_43 sn107_43 11.551961
Rsp106_44 sp106_44 sp107_44 11.551961
Rsn106_44 sn106_44 sn107_44 11.551961
Rsp106_45 sp106_45 sp107_45 11.551961
Rsn106_45 sn106_45 sn107_45 11.551961
Rsp106_46 sp106_46 sp107_46 11.551961
Rsn106_46 sn106_46 sn107_46 11.551961
Rsp106_47 sp106_47 sp107_47 11.551961
Rsn106_47 sn106_47 sn107_47 11.551961
Rsp106_48 sp106_48 sp107_48 11.551961
Rsn106_48 sn106_48 sn107_48 11.551961
Rsp106_49 sp106_49 sp107_49 11.551961
Rsn106_49 sn106_49 sn107_49 11.551961
Rsp106_50 sp106_50 sp107_50 11.551961
Rsn106_50 sn106_50 sn107_50 11.551961
Rsp106_51 sp106_51 sp107_51 11.551961
Rsn106_51 sn106_51 sn107_51 11.551961
Rsp106_52 sp106_52 sp107_52 11.551961
Rsn106_52 sn106_52 sn107_52 11.551961
Rsp106_53 sp106_53 sp107_53 11.551961
Rsn106_53 sn106_53 sn107_53 11.551961
Rsp106_54 sp106_54 sp107_54 11.551961
Rsn106_54 sn106_54 sn107_54 11.551961
Rsp106_55 sp106_55 sp107_55 11.551961
Rsn106_55 sn106_55 sn107_55 11.551961
Rsp106_56 sp106_56 sp107_56 11.551961
Rsn106_56 sn106_56 sn107_56 11.551961
Rsp106_57 sp106_57 sp107_57 11.551961
Rsn106_57 sn106_57 sn107_57 11.551961
Rsp106_58 sp106_58 sp107_58 11.551961
Rsn106_58 sn106_58 sn107_58 11.551961
Rsp106_59 sp106_59 sp107_59 11.551961
Rsn106_59 sn106_59 sn107_59 11.551961
Rsp106_60 sp106_60 sp107_60 11.551961
Rsn106_60 sn106_60 sn107_60 11.551961
Rsp106_61 sp106_61 sp107_61 11.551961
Rsn106_61 sn106_61 sn107_61 11.551961
Rsp106_62 sp106_62 sp107_62 11.551961
Rsn106_62 sn106_62 sn107_62 11.551961
Rsp106_63 sp106_63 sp107_63 11.551961
Rsn106_63 sn106_63 sn107_63 11.551961
Rsp106_64 sp106_64 sp107_64 11.551961
Rsn106_64 sn106_64 sn107_64 11.551961
Rsp106_65 sp106_65 sp107_65 11.551961
Rsn106_65 sn106_65 sn107_65 11.551961
Rsp106_66 sp106_66 sp107_66 11.551961
Rsn106_66 sn106_66 sn107_66 11.551961
Rsp106_67 sp106_67 sp107_67 11.551961
Rsn106_67 sn106_67 sn107_67 11.551961
Rsp106_68 sp106_68 sp107_68 11.551961
Rsn106_68 sn106_68 sn107_68 11.551961
Rsp106_69 sp106_69 sp107_69 11.551961
Rsn106_69 sn106_69 sn107_69 11.551961
Rsp106_70 sp106_70 sp107_70 11.551961
Rsn106_70 sn106_70 sn107_70 11.551961
Rsp106_71 sp106_71 sp107_71 11.551961
Rsn106_71 sn106_71 sn107_71 11.551961
Rsp106_72 sp106_72 sp107_72 11.551961
Rsn106_72 sn106_72 sn107_72 11.551961
Rsp106_73 sp106_73 sp107_73 11.551961
Rsn106_73 sn106_73 sn107_73 11.551961
Rsp106_74 sp106_74 sp107_74 11.551961
Rsn106_74 sn106_74 sn107_74 11.551961
Rsp106_75 sp106_75 sp107_75 11.551961
Rsn106_75 sn106_75 sn107_75 11.551961
Rsp106_76 sp106_76 sp107_76 11.551961
Rsn106_76 sn106_76 sn107_76 11.551961
Rsp106_77 sp106_77 sp107_77 11.551961
Rsn106_77 sn106_77 sn107_77 11.551961
Rsp106_78 sp106_78 sp107_78 11.551961
Rsn106_78 sn106_78 sn107_78 11.551961
Rsp106_79 sp106_79 sp107_79 11.551961
Rsn106_79 sn106_79 sn107_79 11.551961
Rsp106_80 sp106_80 sp107_80 11.551961
Rsn106_80 sn106_80 sn107_80 11.551961
Rsp106_81 sp106_81 sp107_81 11.551961
Rsn106_81 sn106_81 sn107_81 11.551961
Rsp106_82 sp106_82 sp107_82 11.551961
Rsn106_82 sn106_82 sn107_82 11.551961
Rsp106_83 sp106_83 sp107_83 11.551961
Rsn106_83 sn106_83 sn107_83 11.551961
Rsp106_84 sp106_84 sp107_84 11.551961
Rsn106_84 sn106_84 sn107_84 11.551961
Rsp107_1 sp107_1 sp108_1 11.551961
Rsn107_1 sn107_1 sn108_1 11.551961
Rsp107_2 sp107_2 sp108_2 11.551961
Rsn107_2 sn107_2 sn108_2 11.551961
Rsp107_3 sp107_3 sp108_3 11.551961
Rsn107_3 sn107_3 sn108_3 11.551961
Rsp107_4 sp107_4 sp108_4 11.551961
Rsn107_4 sn107_4 sn108_4 11.551961
Rsp107_5 sp107_5 sp108_5 11.551961
Rsn107_5 sn107_5 sn108_5 11.551961
Rsp107_6 sp107_6 sp108_6 11.551961
Rsn107_6 sn107_6 sn108_6 11.551961
Rsp107_7 sp107_7 sp108_7 11.551961
Rsn107_7 sn107_7 sn108_7 11.551961
Rsp107_8 sp107_8 sp108_8 11.551961
Rsn107_8 sn107_8 sn108_8 11.551961
Rsp107_9 sp107_9 sp108_9 11.551961
Rsn107_9 sn107_9 sn108_9 11.551961
Rsp107_10 sp107_10 sp108_10 11.551961
Rsn107_10 sn107_10 sn108_10 11.551961
Rsp107_11 sp107_11 sp108_11 11.551961
Rsn107_11 sn107_11 sn108_11 11.551961
Rsp107_12 sp107_12 sp108_12 11.551961
Rsn107_12 sn107_12 sn108_12 11.551961
Rsp107_13 sp107_13 sp108_13 11.551961
Rsn107_13 sn107_13 sn108_13 11.551961
Rsp107_14 sp107_14 sp108_14 11.551961
Rsn107_14 sn107_14 sn108_14 11.551961
Rsp107_15 sp107_15 sp108_15 11.551961
Rsn107_15 sn107_15 sn108_15 11.551961
Rsp107_16 sp107_16 sp108_16 11.551961
Rsn107_16 sn107_16 sn108_16 11.551961
Rsp107_17 sp107_17 sp108_17 11.551961
Rsn107_17 sn107_17 sn108_17 11.551961
Rsp107_18 sp107_18 sp108_18 11.551961
Rsn107_18 sn107_18 sn108_18 11.551961
Rsp107_19 sp107_19 sp108_19 11.551961
Rsn107_19 sn107_19 sn108_19 11.551961
Rsp107_20 sp107_20 sp108_20 11.551961
Rsn107_20 sn107_20 sn108_20 11.551961
Rsp107_21 sp107_21 sp108_21 11.551961
Rsn107_21 sn107_21 sn108_21 11.551961
Rsp107_22 sp107_22 sp108_22 11.551961
Rsn107_22 sn107_22 sn108_22 11.551961
Rsp107_23 sp107_23 sp108_23 11.551961
Rsn107_23 sn107_23 sn108_23 11.551961
Rsp107_24 sp107_24 sp108_24 11.551961
Rsn107_24 sn107_24 sn108_24 11.551961
Rsp107_25 sp107_25 sp108_25 11.551961
Rsn107_25 sn107_25 sn108_25 11.551961
Rsp107_26 sp107_26 sp108_26 11.551961
Rsn107_26 sn107_26 sn108_26 11.551961
Rsp107_27 sp107_27 sp108_27 11.551961
Rsn107_27 sn107_27 sn108_27 11.551961
Rsp107_28 sp107_28 sp108_28 11.551961
Rsn107_28 sn107_28 sn108_28 11.551961
Rsp107_29 sp107_29 sp108_29 11.551961
Rsn107_29 sn107_29 sn108_29 11.551961
Rsp107_30 sp107_30 sp108_30 11.551961
Rsn107_30 sn107_30 sn108_30 11.551961
Rsp107_31 sp107_31 sp108_31 11.551961
Rsn107_31 sn107_31 sn108_31 11.551961
Rsp107_32 sp107_32 sp108_32 11.551961
Rsn107_32 sn107_32 sn108_32 11.551961
Rsp107_33 sp107_33 sp108_33 11.551961
Rsn107_33 sn107_33 sn108_33 11.551961
Rsp107_34 sp107_34 sp108_34 11.551961
Rsn107_34 sn107_34 sn108_34 11.551961
Rsp107_35 sp107_35 sp108_35 11.551961
Rsn107_35 sn107_35 sn108_35 11.551961
Rsp107_36 sp107_36 sp108_36 11.551961
Rsn107_36 sn107_36 sn108_36 11.551961
Rsp107_37 sp107_37 sp108_37 11.551961
Rsn107_37 sn107_37 sn108_37 11.551961
Rsp107_38 sp107_38 sp108_38 11.551961
Rsn107_38 sn107_38 sn108_38 11.551961
Rsp107_39 sp107_39 sp108_39 11.551961
Rsn107_39 sn107_39 sn108_39 11.551961
Rsp107_40 sp107_40 sp108_40 11.551961
Rsn107_40 sn107_40 sn108_40 11.551961
Rsp107_41 sp107_41 sp108_41 11.551961
Rsn107_41 sn107_41 sn108_41 11.551961
Rsp107_42 sp107_42 sp108_42 11.551961
Rsn107_42 sn107_42 sn108_42 11.551961
Rsp107_43 sp107_43 sp108_43 11.551961
Rsn107_43 sn107_43 sn108_43 11.551961
Rsp107_44 sp107_44 sp108_44 11.551961
Rsn107_44 sn107_44 sn108_44 11.551961
Rsp107_45 sp107_45 sp108_45 11.551961
Rsn107_45 sn107_45 sn108_45 11.551961
Rsp107_46 sp107_46 sp108_46 11.551961
Rsn107_46 sn107_46 sn108_46 11.551961
Rsp107_47 sp107_47 sp108_47 11.551961
Rsn107_47 sn107_47 sn108_47 11.551961
Rsp107_48 sp107_48 sp108_48 11.551961
Rsn107_48 sn107_48 sn108_48 11.551961
Rsp107_49 sp107_49 sp108_49 11.551961
Rsn107_49 sn107_49 sn108_49 11.551961
Rsp107_50 sp107_50 sp108_50 11.551961
Rsn107_50 sn107_50 sn108_50 11.551961
Rsp107_51 sp107_51 sp108_51 11.551961
Rsn107_51 sn107_51 sn108_51 11.551961
Rsp107_52 sp107_52 sp108_52 11.551961
Rsn107_52 sn107_52 sn108_52 11.551961
Rsp107_53 sp107_53 sp108_53 11.551961
Rsn107_53 sn107_53 sn108_53 11.551961
Rsp107_54 sp107_54 sp108_54 11.551961
Rsn107_54 sn107_54 sn108_54 11.551961
Rsp107_55 sp107_55 sp108_55 11.551961
Rsn107_55 sn107_55 sn108_55 11.551961
Rsp107_56 sp107_56 sp108_56 11.551961
Rsn107_56 sn107_56 sn108_56 11.551961
Rsp107_57 sp107_57 sp108_57 11.551961
Rsn107_57 sn107_57 sn108_57 11.551961
Rsp107_58 sp107_58 sp108_58 11.551961
Rsn107_58 sn107_58 sn108_58 11.551961
Rsp107_59 sp107_59 sp108_59 11.551961
Rsn107_59 sn107_59 sn108_59 11.551961
Rsp107_60 sp107_60 sp108_60 11.551961
Rsn107_60 sn107_60 sn108_60 11.551961
Rsp107_61 sp107_61 sp108_61 11.551961
Rsn107_61 sn107_61 sn108_61 11.551961
Rsp107_62 sp107_62 sp108_62 11.551961
Rsn107_62 sn107_62 sn108_62 11.551961
Rsp107_63 sp107_63 sp108_63 11.551961
Rsn107_63 sn107_63 sn108_63 11.551961
Rsp107_64 sp107_64 sp108_64 11.551961
Rsn107_64 sn107_64 sn108_64 11.551961
Rsp107_65 sp107_65 sp108_65 11.551961
Rsn107_65 sn107_65 sn108_65 11.551961
Rsp107_66 sp107_66 sp108_66 11.551961
Rsn107_66 sn107_66 sn108_66 11.551961
Rsp107_67 sp107_67 sp108_67 11.551961
Rsn107_67 sn107_67 sn108_67 11.551961
Rsp107_68 sp107_68 sp108_68 11.551961
Rsn107_68 sn107_68 sn108_68 11.551961
Rsp107_69 sp107_69 sp108_69 11.551961
Rsn107_69 sn107_69 sn108_69 11.551961
Rsp107_70 sp107_70 sp108_70 11.551961
Rsn107_70 sn107_70 sn108_70 11.551961
Rsp107_71 sp107_71 sp108_71 11.551961
Rsn107_71 sn107_71 sn108_71 11.551961
Rsp107_72 sp107_72 sp108_72 11.551961
Rsn107_72 sn107_72 sn108_72 11.551961
Rsp107_73 sp107_73 sp108_73 11.551961
Rsn107_73 sn107_73 sn108_73 11.551961
Rsp107_74 sp107_74 sp108_74 11.551961
Rsn107_74 sn107_74 sn108_74 11.551961
Rsp107_75 sp107_75 sp108_75 11.551961
Rsn107_75 sn107_75 sn108_75 11.551961
Rsp107_76 sp107_76 sp108_76 11.551961
Rsn107_76 sn107_76 sn108_76 11.551961
Rsp107_77 sp107_77 sp108_77 11.551961
Rsn107_77 sn107_77 sn108_77 11.551961
Rsp107_78 sp107_78 sp108_78 11.551961
Rsn107_78 sn107_78 sn108_78 11.551961
Rsp107_79 sp107_79 sp108_79 11.551961
Rsn107_79 sn107_79 sn108_79 11.551961
Rsp107_80 sp107_80 sp108_80 11.551961
Rsn107_80 sn107_80 sn108_80 11.551961
Rsp107_81 sp107_81 sp108_81 11.551961
Rsn107_81 sn107_81 sn108_81 11.551961
Rsp107_82 sp107_82 sp108_82 11.551961
Rsn107_82 sn107_82 sn108_82 11.551961
Rsp107_83 sp107_83 sp108_83 11.551961
Rsn107_83 sn107_83 sn108_83 11.551961
Rsp107_84 sp107_84 sp108_84 11.551961
Rsn107_84 sn107_84 sn108_84 11.551961
Rsp108_1 sp108_1 sp109_1 11.551961
Rsn108_1 sn108_1 sn109_1 11.551961
Rsp108_2 sp108_2 sp109_2 11.551961
Rsn108_2 sn108_2 sn109_2 11.551961
Rsp108_3 sp108_3 sp109_3 11.551961
Rsn108_3 sn108_3 sn109_3 11.551961
Rsp108_4 sp108_4 sp109_4 11.551961
Rsn108_4 sn108_4 sn109_4 11.551961
Rsp108_5 sp108_5 sp109_5 11.551961
Rsn108_5 sn108_5 sn109_5 11.551961
Rsp108_6 sp108_6 sp109_6 11.551961
Rsn108_6 sn108_6 sn109_6 11.551961
Rsp108_7 sp108_7 sp109_7 11.551961
Rsn108_7 sn108_7 sn109_7 11.551961
Rsp108_8 sp108_8 sp109_8 11.551961
Rsn108_8 sn108_8 sn109_8 11.551961
Rsp108_9 sp108_9 sp109_9 11.551961
Rsn108_9 sn108_9 sn109_9 11.551961
Rsp108_10 sp108_10 sp109_10 11.551961
Rsn108_10 sn108_10 sn109_10 11.551961
Rsp108_11 sp108_11 sp109_11 11.551961
Rsn108_11 sn108_11 sn109_11 11.551961
Rsp108_12 sp108_12 sp109_12 11.551961
Rsn108_12 sn108_12 sn109_12 11.551961
Rsp108_13 sp108_13 sp109_13 11.551961
Rsn108_13 sn108_13 sn109_13 11.551961
Rsp108_14 sp108_14 sp109_14 11.551961
Rsn108_14 sn108_14 sn109_14 11.551961
Rsp108_15 sp108_15 sp109_15 11.551961
Rsn108_15 sn108_15 sn109_15 11.551961
Rsp108_16 sp108_16 sp109_16 11.551961
Rsn108_16 sn108_16 sn109_16 11.551961
Rsp108_17 sp108_17 sp109_17 11.551961
Rsn108_17 sn108_17 sn109_17 11.551961
Rsp108_18 sp108_18 sp109_18 11.551961
Rsn108_18 sn108_18 sn109_18 11.551961
Rsp108_19 sp108_19 sp109_19 11.551961
Rsn108_19 sn108_19 sn109_19 11.551961
Rsp108_20 sp108_20 sp109_20 11.551961
Rsn108_20 sn108_20 sn109_20 11.551961
Rsp108_21 sp108_21 sp109_21 11.551961
Rsn108_21 sn108_21 sn109_21 11.551961
Rsp108_22 sp108_22 sp109_22 11.551961
Rsn108_22 sn108_22 sn109_22 11.551961
Rsp108_23 sp108_23 sp109_23 11.551961
Rsn108_23 sn108_23 sn109_23 11.551961
Rsp108_24 sp108_24 sp109_24 11.551961
Rsn108_24 sn108_24 sn109_24 11.551961
Rsp108_25 sp108_25 sp109_25 11.551961
Rsn108_25 sn108_25 sn109_25 11.551961
Rsp108_26 sp108_26 sp109_26 11.551961
Rsn108_26 sn108_26 sn109_26 11.551961
Rsp108_27 sp108_27 sp109_27 11.551961
Rsn108_27 sn108_27 sn109_27 11.551961
Rsp108_28 sp108_28 sp109_28 11.551961
Rsn108_28 sn108_28 sn109_28 11.551961
Rsp108_29 sp108_29 sp109_29 11.551961
Rsn108_29 sn108_29 sn109_29 11.551961
Rsp108_30 sp108_30 sp109_30 11.551961
Rsn108_30 sn108_30 sn109_30 11.551961
Rsp108_31 sp108_31 sp109_31 11.551961
Rsn108_31 sn108_31 sn109_31 11.551961
Rsp108_32 sp108_32 sp109_32 11.551961
Rsn108_32 sn108_32 sn109_32 11.551961
Rsp108_33 sp108_33 sp109_33 11.551961
Rsn108_33 sn108_33 sn109_33 11.551961
Rsp108_34 sp108_34 sp109_34 11.551961
Rsn108_34 sn108_34 sn109_34 11.551961
Rsp108_35 sp108_35 sp109_35 11.551961
Rsn108_35 sn108_35 sn109_35 11.551961
Rsp108_36 sp108_36 sp109_36 11.551961
Rsn108_36 sn108_36 sn109_36 11.551961
Rsp108_37 sp108_37 sp109_37 11.551961
Rsn108_37 sn108_37 sn109_37 11.551961
Rsp108_38 sp108_38 sp109_38 11.551961
Rsn108_38 sn108_38 sn109_38 11.551961
Rsp108_39 sp108_39 sp109_39 11.551961
Rsn108_39 sn108_39 sn109_39 11.551961
Rsp108_40 sp108_40 sp109_40 11.551961
Rsn108_40 sn108_40 sn109_40 11.551961
Rsp108_41 sp108_41 sp109_41 11.551961
Rsn108_41 sn108_41 sn109_41 11.551961
Rsp108_42 sp108_42 sp109_42 11.551961
Rsn108_42 sn108_42 sn109_42 11.551961
Rsp108_43 sp108_43 sp109_43 11.551961
Rsn108_43 sn108_43 sn109_43 11.551961
Rsp108_44 sp108_44 sp109_44 11.551961
Rsn108_44 sn108_44 sn109_44 11.551961
Rsp108_45 sp108_45 sp109_45 11.551961
Rsn108_45 sn108_45 sn109_45 11.551961
Rsp108_46 sp108_46 sp109_46 11.551961
Rsn108_46 sn108_46 sn109_46 11.551961
Rsp108_47 sp108_47 sp109_47 11.551961
Rsn108_47 sn108_47 sn109_47 11.551961
Rsp108_48 sp108_48 sp109_48 11.551961
Rsn108_48 sn108_48 sn109_48 11.551961
Rsp108_49 sp108_49 sp109_49 11.551961
Rsn108_49 sn108_49 sn109_49 11.551961
Rsp108_50 sp108_50 sp109_50 11.551961
Rsn108_50 sn108_50 sn109_50 11.551961
Rsp108_51 sp108_51 sp109_51 11.551961
Rsn108_51 sn108_51 sn109_51 11.551961
Rsp108_52 sp108_52 sp109_52 11.551961
Rsn108_52 sn108_52 sn109_52 11.551961
Rsp108_53 sp108_53 sp109_53 11.551961
Rsn108_53 sn108_53 sn109_53 11.551961
Rsp108_54 sp108_54 sp109_54 11.551961
Rsn108_54 sn108_54 sn109_54 11.551961
Rsp108_55 sp108_55 sp109_55 11.551961
Rsn108_55 sn108_55 sn109_55 11.551961
Rsp108_56 sp108_56 sp109_56 11.551961
Rsn108_56 sn108_56 sn109_56 11.551961
Rsp108_57 sp108_57 sp109_57 11.551961
Rsn108_57 sn108_57 sn109_57 11.551961
Rsp108_58 sp108_58 sp109_58 11.551961
Rsn108_58 sn108_58 sn109_58 11.551961
Rsp108_59 sp108_59 sp109_59 11.551961
Rsn108_59 sn108_59 sn109_59 11.551961
Rsp108_60 sp108_60 sp109_60 11.551961
Rsn108_60 sn108_60 sn109_60 11.551961
Rsp108_61 sp108_61 sp109_61 11.551961
Rsn108_61 sn108_61 sn109_61 11.551961
Rsp108_62 sp108_62 sp109_62 11.551961
Rsn108_62 sn108_62 sn109_62 11.551961
Rsp108_63 sp108_63 sp109_63 11.551961
Rsn108_63 sn108_63 sn109_63 11.551961
Rsp108_64 sp108_64 sp109_64 11.551961
Rsn108_64 sn108_64 sn109_64 11.551961
Rsp108_65 sp108_65 sp109_65 11.551961
Rsn108_65 sn108_65 sn109_65 11.551961
Rsp108_66 sp108_66 sp109_66 11.551961
Rsn108_66 sn108_66 sn109_66 11.551961
Rsp108_67 sp108_67 sp109_67 11.551961
Rsn108_67 sn108_67 sn109_67 11.551961
Rsp108_68 sp108_68 sp109_68 11.551961
Rsn108_68 sn108_68 sn109_68 11.551961
Rsp108_69 sp108_69 sp109_69 11.551961
Rsn108_69 sn108_69 sn109_69 11.551961
Rsp108_70 sp108_70 sp109_70 11.551961
Rsn108_70 sn108_70 sn109_70 11.551961
Rsp108_71 sp108_71 sp109_71 11.551961
Rsn108_71 sn108_71 sn109_71 11.551961
Rsp108_72 sp108_72 sp109_72 11.551961
Rsn108_72 sn108_72 sn109_72 11.551961
Rsp108_73 sp108_73 sp109_73 11.551961
Rsn108_73 sn108_73 sn109_73 11.551961
Rsp108_74 sp108_74 sp109_74 11.551961
Rsn108_74 sn108_74 sn109_74 11.551961
Rsp108_75 sp108_75 sp109_75 11.551961
Rsn108_75 sn108_75 sn109_75 11.551961
Rsp108_76 sp108_76 sp109_76 11.551961
Rsn108_76 sn108_76 sn109_76 11.551961
Rsp108_77 sp108_77 sp109_77 11.551961
Rsn108_77 sn108_77 sn109_77 11.551961
Rsp108_78 sp108_78 sp109_78 11.551961
Rsn108_78 sn108_78 sn109_78 11.551961
Rsp108_79 sp108_79 sp109_79 11.551961
Rsn108_79 sn108_79 sn109_79 11.551961
Rsp108_80 sp108_80 sp109_80 11.551961
Rsn108_80 sn108_80 sn109_80 11.551961
Rsp108_81 sp108_81 sp109_81 11.551961
Rsn108_81 sn108_81 sn109_81 11.551961
Rsp108_82 sp108_82 sp109_82 11.551961
Rsn108_82 sn108_82 sn109_82 11.551961
Rsp108_83 sp108_83 sp109_83 11.551961
Rsn108_83 sn108_83 sn109_83 11.551961
Rsp108_84 sp108_84 sp109_84 11.551961
Rsn108_84 sn108_84 sn109_84 11.551961
Rsp109_1 sp109_1 sp110_1 11.551961
Rsn109_1 sn109_1 sn110_1 11.551961
Rsp109_2 sp109_2 sp110_2 11.551961
Rsn109_2 sn109_2 sn110_2 11.551961
Rsp109_3 sp109_3 sp110_3 11.551961
Rsn109_3 sn109_3 sn110_3 11.551961
Rsp109_4 sp109_4 sp110_4 11.551961
Rsn109_4 sn109_4 sn110_4 11.551961
Rsp109_5 sp109_5 sp110_5 11.551961
Rsn109_5 sn109_5 sn110_5 11.551961
Rsp109_6 sp109_6 sp110_6 11.551961
Rsn109_6 sn109_6 sn110_6 11.551961
Rsp109_7 sp109_7 sp110_7 11.551961
Rsn109_7 sn109_7 sn110_7 11.551961
Rsp109_8 sp109_8 sp110_8 11.551961
Rsn109_8 sn109_8 sn110_8 11.551961
Rsp109_9 sp109_9 sp110_9 11.551961
Rsn109_9 sn109_9 sn110_9 11.551961
Rsp109_10 sp109_10 sp110_10 11.551961
Rsn109_10 sn109_10 sn110_10 11.551961
Rsp109_11 sp109_11 sp110_11 11.551961
Rsn109_11 sn109_11 sn110_11 11.551961
Rsp109_12 sp109_12 sp110_12 11.551961
Rsn109_12 sn109_12 sn110_12 11.551961
Rsp109_13 sp109_13 sp110_13 11.551961
Rsn109_13 sn109_13 sn110_13 11.551961
Rsp109_14 sp109_14 sp110_14 11.551961
Rsn109_14 sn109_14 sn110_14 11.551961
Rsp109_15 sp109_15 sp110_15 11.551961
Rsn109_15 sn109_15 sn110_15 11.551961
Rsp109_16 sp109_16 sp110_16 11.551961
Rsn109_16 sn109_16 sn110_16 11.551961
Rsp109_17 sp109_17 sp110_17 11.551961
Rsn109_17 sn109_17 sn110_17 11.551961
Rsp109_18 sp109_18 sp110_18 11.551961
Rsn109_18 sn109_18 sn110_18 11.551961
Rsp109_19 sp109_19 sp110_19 11.551961
Rsn109_19 sn109_19 sn110_19 11.551961
Rsp109_20 sp109_20 sp110_20 11.551961
Rsn109_20 sn109_20 sn110_20 11.551961
Rsp109_21 sp109_21 sp110_21 11.551961
Rsn109_21 sn109_21 sn110_21 11.551961
Rsp109_22 sp109_22 sp110_22 11.551961
Rsn109_22 sn109_22 sn110_22 11.551961
Rsp109_23 sp109_23 sp110_23 11.551961
Rsn109_23 sn109_23 sn110_23 11.551961
Rsp109_24 sp109_24 sp110_24 11.551961
Rsn109_24 sn109_24 sn110_24 11.551961
Rsp109_25 sp109_25 sp110_25 11.551961
Rsn109_25 sn109_25 sn110_25 11.551961
Rsp109_26 sp109_26 sp110_26 11.551961
Rsn109_26 sn109_26 sn110_26 11.551961
Rsp109_27 sp109_27 sp110_27 11.551961
Rsn109_27 sn109_27 sn110_27 11.551961
Rsp109_28 sp109_28 sp110_28 11.551961
Rsn109_28 sn109_28 sn110_28 11.551961
Rsp109_29 sp109_29 sp110_29 11.551961
Rsn109_29 sn109_29 sn110_29 11.551961
Rsp109_30 sp109_30 sp110_30 11.551961
Rsn109_30 sn109_30 sn110_30 11.551961
Rsp109_31 sp109_31 sp110_31 11.551961
Rsn109_31 sn109_31 sn110_31 11.551961
Rsp109_32 sp109_32 sp110_32 11.551961
Rsn109_32 sn109_32 sn110_32 11.551961
Rsp109_33 sp109_33 sp110_33 11.551961
Rsn109_33 sn109_33 sn110_33 11.551961
Rsp109_34 sp109_34 sp110_34 11.551961
Rsn109_34 sn109_34 sn110_34 11.551961
Rsp109_35 sp109_35 sp110_35 11.551961
Rsn109_35 sn109_35 sn110_35 11.551961
Rsp109_36 sp109_36 sp110_36 11.551961
Rsn109_36 sn109_36 sn110_36 11.551961
Rsp109_37 sp109_37 sp110_37 11.551961
Rsn109_37 sn109_37 sn110_37 11.551961
Rsp109_38 sp109_38 sp110_38 11.551961
Rsn109_38 sn109_38 sn110_38 11.551961
Rsp109_39 sp109_39 sp110_39 11.551961
Rsn109_39 sn109_39 sn110_39 11.551961
Rsp109_40 sp109_40 sp110_40 11.551961
Rsn109_40 sn109_40 sn110_40 11.551961
Rsp109_41 sp109_41 sp110_41 11.551961
Rsn109_41 sn109_41 sn110_41 11.551961
Rsp109_42 sp109_42 sp110_42 11.551961
Rsn109_42 sn109_42 sn110_42 11.551961
Rsp109_43 sp109_43 sp110_43 11.551961
Rsn109_43 sn109_43 sn110_43 11.551961
Rsp109_44 sp109_44 sp110_44 11.551961
Rsn109_44 sn109_44 sn110_44 11.551961
Rsp109_45 sp109_45 sp110_45 11.551961
Rsn109_45 sn109_45 sn110_45 11.551961
Rsp109_46 sp109_46 sp110_46 11.551961
Rsn109_46 sn109_46 sn110_46 11.551961
Rsp109_47 sp109_47 sp110_47 11.551961
Rsn109_47 sn109_47 sn110_47 11.551961
Rsp109_48 sp109_48 sp110_48 11.551961
Rsn109_48 sn109_48 sn110_48 11.551961
Rsp109_49 sp109_49 sp110_49 11.551961
Rsn109_49 sn109_49 sn110_49 11.551961
Rsp109_50 sp109_50 sp110_50 11.551961
Rsn109_50 sn109_50 sn110_50 11.551961
Rsp109_51 sp109_51 sp110_51 11.551961
Rsn109_51 sn109_51 sn110_51 11.551961
Rsp109_52 sp109_52 sp110_52 11.551961
Rsn109_52 sn109_52 sn110_52 11.551961
Rsp109_53 sp109_53 sp110_53 11.551961
Rsn109_53 sn109_53 sn110_53 11.551961
Rsp109_54 sp109_54 sp110_54 11.551961
Rsn109_54 sn109_54 sn110_54 11.551961
Rsp109_55 sp109_55 sp110_55 11.551961
Rsn109_55 sn109_55 sn110_55 11.551961
Rsp109_56 sp109_56 sp110_56 11.551961
Rsn109_56 sn109_56 sn110_56 11.551961
Rsp109_57 sp109_57 sp110_57 11.551961
Rsn109_57 sn109_57 sn110_57 11.551961
Rsp109_58 sp109_58 sp110_58 11.551961
Rsn109_58 sn109_58 sn110_58 11.551961
Rsp109_59 sp109_59 sp110_59 11.551961
Rsn109_59 sn109_59 sn110_59 11.551961
Rsp109_60 sp109_60 sp110_60 11.551961
Rsn109_60 sn109_60 sn110_60 11.551961
Rsp109_61 sp109_61 sp110_61 11.551961
Rsn109_61 sn109_61 sn110_61 11.551961
Rsp109_62 sp109_62 sp110_62 11.551961
Rsn109_62 sn109_62 sn110_62 11.551961
Rsp109_63 sp109_63 sp110_63 11.551961
Rsn109_63 sn109_63 sn110_63 11.551961
Rsp109_64 sp109_64 sp110_64 11.551961
Rsn109_64 sn109_64 sn110_64 11.551961
Rsp109_65 sp109_65 sp110_65 11.551961
Rsn109_65 sn109_65 sn110_65 11.551961
Rsp109_66 sp109_66 sp110_66 11.551961
Rsn109_66 sn109_66 sn110_66 11.551961
Rsp109_67 sp109_67 sp110_67 11.551961
Rsn109_67 sn109_67 sn110_67 11.551961
Rsp109_68 sp109_68 sp110_68 11.551961
Rsn109_68 sn109_68 sn110_68 11.551961
Rsp109_69 sp109_69 sp110_69 11.551961
Rsn109_69 sn109_69 sn110_69 11.551961
Rsp109_70 sp109_70 sp110_70 11.551961
Rsn109_70 sn109_70 sn110_70 11.551961
Rsp109_71 sp109_71 sp110_71 11.551961
Rsn109_71 sn109_71 sn110_71 11.551961
Rsp109_72 sp109_72 sp110_72 11.551961
Rsn109_72 sn109_72 sn110_72 11.551961
Rsp109_73 sp109_73 sp110_73 11.551961
Rsn109_73 sn109_73 sn110_73 11.551961
Rsp109_74 sp109_74 sp110_74 11.551961
Rsn109_74 sn109_74 sn110_74 11.551961
Rsp109_75 sp109_75 sp110_75 11.551961
Rsn109_75 sn109_75 sn110_75 11.551961
Rsp109_76 sp109_76 sp110_76 11.551961
Rsn109_76 sn109_76 sn110_76 11.551961
Rsp109_77 sp109_77 sp110_77 11.551961
Rsn109_77 sn109_77 sn110_77 11.551961
Rsp109_78 sp109_78 sp110_78 11.551961
Rsn109_78 sn109_78 sn110_78 11.551961
Rsp109_79 sp109_79 sp110_79 11.551961
Rsn109_79 sn109_79 sn110_79 11.551961
Rsp109_80 sp109_80 sp110_80 11.551961
Rsn109_80 sn109_80 sn110_80 11.551961
Rsp109_81 sp109_81 sp110_81 11.551961
Rsn109_81 sn109_81 sn110_81 11.551961
Rsp109_82 sp109_82 sp110_82 11.551961
Rsn109_82 sn109_82 sn110_82 11.551961
Rsp109_83 sp109_83 sp110_83 11.551961
Rsn109_83 sn109_83 sn110_83 11.551961
Rsp109_84 sp109_84 sp110_84 11.551961
Rsn109_84 sn109_84 sn110_84 11.551961
Rsp110_1 sp110_1 sp111_1 11.551961
Rsn110_1 sn110_1 sn111_1 11.551961
Rsp110_2 sp110_2 sp111_2 11.551961
Rsn110_2 sn110_2 sn111_2 11.551961
Rsp110_3 sp110_3 sp111_3 11.551961
Rsn110_3 sn110_3 sn111_3 11.551961
Rsp110_4 sp110_4 sp111_4 11.551961
Rsn110_4 sn110_4 sn111_4 11.551961
Rsp110_5 sp110_5 sp111_5 11.551961
Rsn110_5 sn110_5 sn111_5 11.551961
Rsp110_6 sp110_6 sp111_6 11.551961
Rsn110_6 sn110_6 sn111_6 11.551961
Rsp110_7 sp110_7 sp111_7 11.551961
Rsn110_7 sn110_7 sn111_7 11.551961
Rsp110_8 sp110_8 sp111_8 11.551961
Rsn110_8 sn110_8 sn111_8 11.551961
Rsp110_9 sp110_9 sp111_9 11.551961
Rsn110_9 sn110_9 sn111_9 11.551961
Rsp110_10 sp110_10 sp111_10 11.551961
Rsn110_10 sn110_10 sn111_10 11.551961
Rsp110_11 sp110_11 sp111_11 11.551961
Rsn110_11 sn110_11 sn111_11 11.551961
Rsp110_12 sp110_12 sp111_12 11.551961
Rsn110_12 sn110_12 sn111_12 11.551961
Rsp110_13 sp110_13 sp111_13 11.551961
Rsn110_13 sn110_13 sn111_13 11.551961
Rsp110_14 sp110_14 sp111_14 11.551961
Rsn110_14 sn110_14 sn111_14 11.551961
Rsp110_15 sp110_15 sp111_15 11.551961
Rsn110_15 sn110_15 sn111_15 11.551961
Rsp110_16 sp110_16 sp111_16 11.551961
Rsn110_16 sn110_16 sn111_16 11.551961
Rsp110_17 sp110_17 sp111_17 11.551961
Rsn110_17 sn110_17 sn111_17 11.551961
Rsp110_18 sp110_18 sp111_18 11.551961
Rsn110_18 sn110_18 sn111_18 11.551961
Rsp110_19 sp110_19 sp111_19 11.551961
Rsn110_19 sn110_19 sn111_19 11.551961
Rsp110_20 sp110_20 sp111_20 11.551961
Rsn110_20 sn110_20 sn111_20 11.551961
Rsp110_21 sp110_21 sp111_21 11.551961
Rsn110_21 sn110_21 sn111_21 11.551961
Rsp110_22 sp110_22 sp111_22 11.551961
Rsn110_22 sn110_22 sn111_22 11.551961
Rsp110_23 sp110_23 sp111_23 11.551961
Rsn110_23 sn110_23 sn111_23 11.551961
Rsp110_24 sp110_24 sp111_24 11.551961
Rsn110_24 sn110_24 sn111_24 11.551961
Rsp110_25 sp110_25 sp111_25 11.551961
Rsn110_25 sn110_25 sn111_25 11.551961
Rsp110_26 sp110_26 sp111_26 11.551961
Rsn110_26 sn110_26 sn111_26 11.551961
Rsp110_27 sp110_27 sp111_27 11.551961
Rsn110_27 sn110_27 sn111_27 11.551961
Rsp110_28 sp110_28 sp111_28 11.551961
Rsn110_28 sn110_28 sn111_28 11.551961
Rsp110_29 sp110_29 sp111_29 11.551961
Rsn110_29 sn110_29 sn111_29 11.551961
Rsp110_30 sp110_30 sp111_30 11.551961
Rsn110_30 sn110_30 sn111_30 11.551961
Rsp110_31 sp110_31 sp111_31 11.551961
Rsn110_31 sn110_31 sn111_31 11.551961
Rsp110_32 sp110_32 sp111_32 11.551961
Rsn110_32 sn110_32 sn111_32 11.551961
Rsp110_33 sp110_33 sp111_33 11.551961
Rsn110_33 sn110_33 sn111_33 11.551961
Rsp110_34 sp110_34 sp111_34 11.551961
Rsn110_34 sn110_34 sn111_34 11.551961
Rsp110_35 sp110_35 sp111_35 11.551961
Rsn110_35 sn110_35 sn111_35 11.551961
Rsp110_36 sp110_36 sp111_36 11.551961
Rsn110_36 sn110_36 sn111_36 11.551961
Rsp110_37 sp110_37 sp111_37 11.551961
Rsn110_37 sn110_37 sn111_37 11.551961
Rsp110_38 sp110_38 sp111_38 11.551961
Rsn110_38 sn110_38 sn111_38 11.551961
Rsp110_39 sp110_39 sp111_39 11.551961
Rsn110_39 sn110_39 sn111_39 11.551961
Rsp110_40 sp110_40 sp111_40 11.551961
Rsn110_40 sn110_40 sn111_40 11.551961
Rsp110_41 sp110_41 sp111_41 11.551961
Rsn110_41 sn110_41 sn111_41 11.551961
Rsp110_42 sp110_42 sp111_42 11.551961
Rsn110_42 sn110_42 sn111_42 11.551961
Rsp110_43 sp110_43 sp111_43 11.551961
Rsn110_43 sn110_43 sn111_43 11.551961
Rsp110_44 sp110_44 sp111_44 11.551961
Rsn110_44 sn110_44 sn111_44 11.551961
Rsp110_45 sp110_45 sp111_45 11.551961
Rsn110_45 sn110_45 sn111_45 11.551961
Rsp110_46 sp110_46 sp111_46 11.551961
Rsn110_46 sn110_46 sn111_46 11.551961
Rsp110_47 sp110_47 sp111_47 11.551961
Rsn110_47 sn110_47 sn111_47 11.551961
Rsp110_48 sp110_48 sp111_48 11.551961
Rsn110_48 sn110_48 sn111_48 11.551961
Rsp110_49 sp110_49 sp111_49 11.551961
Rsn110_49 sn110_49 sn111_49 11.551961
Rsp110_50 sp110_50 sp111_50 11.551961
Rsn110_50 sn110_50 sn111_50 11.551961
Rsp110_51 sp110_51 sp111_51 11.551961
Rsn110_51 sn110_51 sn111_51 11.551961
Rsp110_52 sp110_52 sp111_52 11.551961
Rsn110_52 sn110_52 sn111_52 11.551961
Rsp110_53 sp110_53 sp111_53 11.551961
Rsn110_53 sn110_53 sn111_53 11.551961
Rsp110_54 sp110_54 sp111_54 11.551961
Rsn110_54 sn110_54 sn111_54 11.551961
Rsp110_55 sp110_55 sp111_55 11.551961
Rsn110_55 sn110_55 sn111_55 11.551961
Rsp110_56 sp110_56 sp111_56 11.551961
Rsn110_56 sn110_56 sn111_56 11.551961
Rsp110_57 sp110_57 sp111_57 11.551961
Rsn110_57 sn110_57 sn111_57 11.551961
Rsp110_58 sp110_58 sp111_58 11.551961
Rsn110_58 sn110_58 sn111_58 11.551961
Rsp110_59 sp110_59 sp111_59 11.551961
Rsn110_59 sn110_59 sn111_59 11.551961
Rsp110_60 sp110_60 sp111_60 11.551961
Rsn110_60 sn110_60 sn111_60 11.551961
Rsp110_61 sp110_61 sp111_61 11.551961
Rsn110_61 sn110_61 sn111_61 11.551961
Rsp110_62 sp110_62 sp111_62 11.551961
Rsn110_62 sn110_62 sn111_62 11.551961
Rsp110_63 sp110_63 sp111_63 11.551961
Rsn110_63 sn110_63 sn111_63 11.551961
Rsp110_64 sp110_64 sp111_64 11.551961
Rsn110_64 sn110_64 sn111_64 11.551961
Rsp110_65 sp110_65 sp111_65 11.551961
Rsn110_65 sn110_65 sn111_65 11.551961
Rsp110_66 sp110_66 sp111_66 11.551961
Rsn110_66 sn110_66 sn111_66 11.551961
Rsp110_67 sp110_67 sp111_67 11.551961
Rsn110_67 sn110_67 sn111_67 11.551961
Rsp110_68 sp110_68 sp111_68 11.551961
Rsn110_68 sn110_68 sn111_68 11.551961
Rsp110_69 sp110_69 sp111_69 11.551961
Rsn110_69 sn110_69 sn111_69 11.551961
Rsp110_70 sp110_70 sp111_70 11.551961
Rsn110_70 sn110_70 sn111_70 11.551961
Rsp110_71 sp110_71 sp111_71 11.551961
Rsn110_71 sn110_71 sn111_71 11.551961
Rsp110_72 sp110_72 sp111_72 11.551961
Rsn110_72 sn110_72 sn111_72 11.551961
Rsp110_73 sp110_73 sp111_73 11.551961
Rsn110_73 sn110_73 sn111_73 11.551961
Rsp110_74 sp110_74 sp111_74 11.551961
Rsn110_74 sn110_74 sn111_74 11.551961
Rsp110_75 sp110_75 sp111_75 11.551961
Rsn110_75 sn110_75 sn111_75 11.551961
Rsp110_76 sp110_76 sp111_76 11.551961
Rsn110_76 sn110_76 sn111_76 11.551961
Rsp110_77 sp110_77 sp111_77 11.551961
Rsn110_77 sn110_77 sn111_77 11.551961
Rsp110_78 sp110_78 sp111_78 11.551961
Rsn110_78 sn110_78 sn111_78 11.551961
Rsp110_79 sp110_79 sp111_79 11.551961
Rsn110_79 sn110_79 sn111_79 11.551961
Rsp110_80 sp110_80 sp111_80 11.551961
Rsn110_80 sn110_80 sn111_80 11.551961
Rsp110_81 sp110_81 sp111_81 11.551961
Rsn110_81 sn110_81 sn111_81 11.551961
Rsp110_82 sp110_82 sp111_82 11.551961
Rsn110_82 sn110_82 sn111_82 11.551961
Rsp110_83 sp110_83 sp111_83 11.551961
Rsn110_83 sn110_83 sn111_83 11.551961
Rsp110_84 sp110_84 sp111_84 11.551961
Rsn110_84 sn110_84 sn111_84 11.551961
Rsp111_1 sp111_1 sp112_1 11.551961
Rsn111_1 sn111_1 sn112_1 11.551961
Rsp111_2 sp111_2 sp112_2 11.551961
Rsn111_2 sn111_2 sn112_2 11.551961
Rsp111_3 sp111_3 sp112_3 11.551961
Rsn111_3 sn111_3 sn112_3 11.551961
Rsp111_4 sp111_4 sp112_4 11.551961
Rsn111_4 sn111_4 sn112_4 11.551961
Rsp111_5 sp111_5 sp112_5 11.551961
Rsn111_5 sn111_5 sn112_5 11.551961
Rsp111_6 sp111_6 sp112_6 11.551961
Rsn111_6 sn111_6 sn112_6 11.551961
Rsp111_7 sp111_7 sp112_7 11.551961
Rsn111_7 sn111_7 sn112_7 11.551961
Rsp111_8 sp111_8 sp112_8 11.551961
Rsn111_8 sn111_8 sn112_8 11.551961
Rsp111_9 sp111_9 sp112_9 11.551961
Rsn111_9 sn111_9 sn112_9 11.551961
Rsp111_10 sp111_10 sp112_10 11.551961
Rsn111_10 sn111_10 sn112_10 11.551961
Rsp111_11 sp111_11 sp112_11 11.551961
Rsn111_11 sn111_11 sn112_11 11.551961
Rsp111_12 sp111_12 sp112_12 11.551961
Rsn111_12 sn111_12 sn112_12 11.551961
Rsp111_13 sp111_13 sp112_13 11.551961
Rsn111_13 sn111_13 sn112_13 11.551961
Rsp111_14 sp111_14 sp112_14 11.551961
Rsn111_14 sn111_14 sn112_14 11.551961
Rsp111_15 sp111_15 sp112_15 11.551961
Rsn111_15 sn111_15 sn112_15 11.551961
Rsp111_16 sp111_16 sp112_16 11.551961
Rsn111_16 sn111_16 sn112_16 11.551961
Rsp111_17 sp111_17 sp112_17 11.551961
Rsn111_17 sn111_17 sn112_17 11.551961
Rsp111_18 sp111_18 sp112_18 11.551961
Rsn111_18 sn111_18 sn112_18 11.551961
Rsp111_19 sp111_19 sp112_19 11.551961
Rsn111_19 sn111_19 sn112_19 11.551961
Rsp111_20 sp111_20 sp112_20 11.551961
Rsn111_20 sn111_20 sn112_20 11.551961
Rsp111_21 sp111_21 sp112_21 11.551961
Rsn111_21 sn111_21 sn112_21 11.551961
Rsp111_22 sp111_22 sp112_22 11.551961
Rsn111_22 sn111_22 sn112_22 11.551961
Rsp111_23 sp111_23 sp112_23 11.551961
Rsn111_23 sn111_23 sn112_23 11.551961
Rsp111_24 sp111_24 sp112_24 11.551961
Rsn111_24 sn111_24 sn112_24 11.551961
Rsp111_25 sp111_25 sp112_25 11.551961
Rsn111_25 sn111_25 sn112_25 11.551961
Rsp111_26 sp111_26 sp112_26 11.551961
Rsn111_26 sn111_26 sn112_26 11.551961
Rsp111_27 sp111_27 sp112_27 11.551961
Rsn111_27 sn111_27 sn112_27 11.551961
Rsp111_28 sp111_28 sp112_28 11.551961
Rsn111_28 sn111_28 sn112_28 11.551961
Rsp111_29 sp111_29 sp112_29 11.551961
Rsn111_29 sn111_29 sn112_29 11.551961
Rsp111_30 sp111_30 sp112_30 11.551961
Rsn111_30 sn111_30 sn112_30 11.551961
Rsp111_31 sp111_31 sp112_31 11.551961
Rsn111_31 sn111_31 sn112_31 11.551961
Rsp111_32 sp111_32 sp112_32 11.551961
Rsn111_32 sn111_32 sn112_32 11.551961
Rsp111_33 sp111_33 sp112_33 11.551961
Rsn111_33 sn111_33 sn112_33 11.551961
Rsp111_34 sp111_34 sp112_34 11.551961
Rsn111_34 sn111_34 sn112_34 11.551961
Rsp111_35 sp111_35 sp112_35 11.551961
Rsn111_35 sn111_35 sn112_35 11.551961
Rsp111_36 sp111_36 sp112_36 11.551961
Rsn111_36 sn111_36 sn112_36 11.551961
Rsp111_37 sp111_37 sp112_37 11.551961
Rsn111_37 sn111_37 sn112_37 11.551961
Rsp111_38 sp111_38 sp112_38 11.551961
Rsn111_38 sn111_38 sn112_38 11.551961
Rsp111_39 sp111_39 sp112_39 11.551961
Rsn111_39 sn111_39 sn112_39 11.551961
Rsp111_40 sp111_40 sp112_40 11.551961
Rsn111_40 sn111_40 sn112_40 11.551961
Rsp111_41 sp111_41 sp112_41 11.551961
Rsn111_41 sn111_41 sn112_41 11.551961
Rsp111_42 sp111_42 sp112_42 11.551961
Rsn111_42 sn111_42 sn112_42 11.551961
Rsp111_43 sp111_43 sp112_43 11.551961
Rsn111_43 sn111_43 sn112_43 11.551961
Rsp111_44 sp111_44 sp112_44 11.551961
Rsn111_44 sn111_44 sn112_44 11.551961
Rsp111_45 sp111_45 sp112_45 11.551961
Rsn111_45 sn111_45 sn112_45 11.551961
Rsp111_46 sp111_46 sp112_46 11.551961
Rsn111_46 sn111_46 sn112_46 11.551961
Rsp111_47 sp111_47 sp112_47 11.551961
Rsn111_47 sn111_47 sn112_47 11.551961
Rsp111_48 sp111_48 sp112_48 11.551961
Rsn111_48 sn111_48 sn112_48 11.551961
Rsp111_49 sp111_49 sp112_49 11.551961
Rsn111_49 sn111_49 sn112_49 11.551961
Rsp111_50 sp111_50 sp112_50 11.551961
Rsn111_50 sn111_50 sn112_50 11.551961
Rsp111_51 sp111_51 sp112_51 11.551961
Rsn111_51 sn111_51 sn112_51 11.551961
Rsp111_52 sp111_52 sp112_52 11.551961
Rsn111_52 sn111_52 sn112_52 11.551961
Rsp111_53 sp111_53 sp112_53 11.551961
Rsn111_53 sn111_53 sn112_53 11.551961
Rsp111_54 sp111_54 sp112_54 11.551961
Rsn111_54 sn111_54 sn112_54 11.551961
Rsp111_55 sp111_55 sp112_55 11.551961
Rsn111_55 sn111_55 sn112_55 11.551961
Rsp111_56 sp111_56 sp112_56 11.551961
Rsn111_56 sn111_56 sn112_56 11.551961
Rsp111_57 sp111_57 sp112_57 11.551961
Rsn111_57 sn111_57 sn112_57 11.551961
Rsp111_58 sp111_58 sp112_58 11.551961
Rsn111_58 sn111_58 sn112_58 11.551961
Rsp111_59 sp111_59 sp112_59 11.551961
Rsn111_59 sn111_59 sn112_59 11.551961
Rsp111_60 sp111_60 sp112_60 11.551961
Rsn111_60 sn111_60 sn112_60 11.551961
Rsp111_61 sp111_61 sp112_61 11.551961
Rsn111_61 sn111_61 sn112_61 11.551961
Rsp111_62 sp111_62 sp112_62 11.551961
Rsn111_62 sn111_62 sn112_62 11.551961
Rsp111_63 sp111_63 sp112_63 11.551961
Rsn111_63 sn111_63 sn112_63 11.551961
Rsp111_64 sp111_64 sp112_64 11.551961
Rsn111_64 sn111_64 sn112_64 11.551961
Rsp111_65 sp111_65 sp112_65 11.551961
Rsn111_65 sn111_65 sn112_65 11.551961
Rsp111_66 sp111_66 sp112_66 11.551961
Rsn111_66 sn111_66 sn112_66 11.551961
Rsp111_67 sp111_67 sp112_67 11.551961
Rsn111_67 sn111_67 sn112_67 11.551961
Rsp111_68 sp111_68 sp112_68 11.551961
Rsn111_68 sn111_68 sn112_68 11.551961
Rsp111_69 sp111_69 sp112_69 11.551961
Rsn111_69 sn111_69 sn112_69 11.551961
Rsp111_70 sp111_70 sp112_70 11.551961
Rsn111_70 sn111_70 sn112_70 11.551961
Rsp111_71 sp111_71 sp112_71 11.551961
Rsn111_71 sn111_71 sn112_71 11.551961
Rsp111_72 sp111_72 sp112_72 11.551961
Rsn111_72 sn111_72 sn112_72 11.551961
Rsp111_73 sp111_73 sp112_73 11.551961
Rsn111_73 sn111_73 sn112_73 11.551961
Rsp111_74 sp111_74 sp112_74 11.551961
Rsn111_74 sn111_74 sn112_74 11.551961
Rsp111_75 sp111_75 sp112_75 11.551961
Rsn111_75 sn111_75 sn112_75 11.551961
Rsp111_76 sp111_76 sp112_76 11.551961
Rsn111_76 sn111_76 sn112_76 11.551961
Rsp111_77 sp111_77 sp112_77 11.551961
Rsn111_77 sn111_77 sn112_77 11.551961
Rsp111_78 sp111_78 sp112_78 11.551961
Rsn111_78 sn111_78 sn112_78 11.551961
Rsp111_79 sp111_79 sp112_79 11.551961
Rsn111_79 sn111_79 sn112_79 11.551961
Rsp111_80 sp111_80 sp112_80 11.551961
Rsn111_80 sn111_80 sn112_80 11.551961
Rsp111_81 sp111_81 sp112_81 11.551961
Rsn111_81 sn111_81 sn112_81 11.551961
Rsp111_82 sp111_82 sp112_82 11.551961
Rsn111_82 sn111_82 sn112_82 11.551961
Rsp111_83 sp111_83 sp112_83 11.551961
Rsn111_83 sn111_83 sn112_83 11.551961
Rsp111_84 sp111_84 sp112_84 11.551961
Rsn111_84 sn111_84 sn112_84 11.551961
Rsp112_1 sp112_1 sp113_1 11.551961
Rsn112_1 sn112_1 sn113_1 11.551961
Rsp112_2 sp112_2 sp113_2 11.551961
Rsn112_2 sn112_2 sn113_2 11.551961
Rsp112_3 sp112_3 sp113_3 11.551961
Rsn112_3 sn112_3 sn113_3 11.551961
Rsp112_4 sp112_4 sp113_4 11.551961
Rsn112_4 sn112_4 sn113_4 11.551961
Rsp112_5 sp112_5 sp113_5 11.551961
Rsn112_5 sn112_5 sn113_5 11.551961
Rsp112_6 sp112_6 sp113_6 11.551961
Rsn112_6 sn112_6 sn113_6 11.551961
Rsp112_7 sp112_7 sp113_7 11.551961
Rsn112_7 sn112_7 sn113_7 11.551961
Rsp112_8 sp112_8 sp113_8 11.551961
Rsn112_8 sn112_8 sn113_8 11.551961
Rsp112_9 sp112_9 sp113_9 11.551961
Rsn112_9 sn112_9 sn113_9 11.551961
Rsp112_10 sp112_10 sp113_10 11.551961
Rsn112_10 sn112_10 sn113_10 11.551961
Rsp112_11 sp112_11 sp113_11 11.551961
Rsn112_11 sn112_11 sn113_11 11.551961
Rsp112_12 sp112_12 sp113_12 11.551961
Rsn112_12 sn112_12 sn113_12 11.551961
Rsp112_13 sp112_13 sp113_13 11.551961
Rsn112_13 sn112_13 sn113_13 11.551961
Rsp112_14 sp112_14 sp113_14 11.551961
Rsn112_14 sn112_14 sn113_14 11.551961
Rsp112_15 sp112_15 sp113_15 11.551961
Rsn112_15 sn112_15 sn113_15 11.551961
Rsp112_16 sp112_16 sp113_16 11.551961
Rsn112_16 sn112_16 sn113_16 11.551961
Rsp112_17 sp112_17 sp113_17 11.551961
Rsn112_17 sn112_17 sn113_17 11.551961
Rsp112_18 sp112_18 sp113_18 11.551961
Rsn112_18 sn112_18 sn113_18 11.551961
Rsp112_19 sp112_19 sp113_19 11.551961
Rsn112_19 sn112_19 sn113_19 11.551961
Rsp112_20 sp112_20 sp113_20 11.551961
Rsn112_20 sn112_20 sn113_20 11.551961
Rsp112_21 sp112_21 sp113_21 11.551961
Rsn112_21 sn112_21 sn113_21 11.551961
Rsp112_22 sp112_22 sp113_22 11.551961
Rsn112_22 sn112_22 sn113_22 11.551961
Rsp112_23 sp112_23 sp113_23 11.551961
Rsn112_23 sn112_23 sn113_23 11.551961
Rsp112_24 sp112_24 sp113_24 11.551961
Rsn112_24 sn112_24 sn113_24 11.551961
Rsp112_25 sp112_25 sp113_25 11.551961
Rsn112_25 sn112_25 sn113_25 11.551961
Rsp112_26 sp112_26 sp113_26 11.551961
Rsn112_26 sn112_26 sn113_26 11.551961
Rsp112_27 sp112_27 sp113_27 11.551961
Rsn112_27 sn112_27 sn113_27 11.551961
Rsp112_28 sp112_28 sp113_28 11.551961
Rsn112_28 sn112_28 sn113_28 11.551961
Rsp112_29 sp112_29 sp113_29 11.551961
Rsn112_29 sn112_29 sn113_29 11.551961
Rsp112_30 sp112_30 sp113_30 11.551961
Rsn112_30 sn112_30 sn113_30 11.551961
Rsp112_31 sp112_31 sp113_31 11.551961
Rsn112_31 sn112_31 sn113_31 11.551961
Rsp112_32 sp112_32 sp113_32 11.551961
Rsn112_32 sn112_32 sn113_32 11.551961
Rsp112_33 sp112_33 sp113_33 11.551961
Rsn112_33 sn112_33 sn113_33 11.551961
Rsp112_34 sp112_34 sp113_34 11.551961
Rsn112_34 sn112_34 sn113_34 11.551961
Rsp112_35 sp112_35 sp113_35 11.551961
Rsn112_35 sn112_35 sn113_35 11.551961
Rsp112_36 sp112_36 sp113_36 11.551961
Rsn112_36 sn112_36 sn113_36 11.551961
Rsp112_37 sp112_37 sp113_37 11.551961
Rsn112_37 sn112_37 sn113_37 11.551961
Rsp112_38 sp112_38 sp113_38 11.551961
Rsn112_38 sn112_38 sn113_38 11.551961
Rsp112_39 sp112_39 sp113_39 11.551961
Rsn112_39 sn112_39 sn113_39 11.551961
Rsp112_40 sp112_40 sp113_40 11.551961
Rsn112_40 sn112_40 sn113_40 11.551961
Rsp112_41 sp112_41 sp113_41 11.551961
Rsn112_41 sn112_41 sn113_41 11.551961
Rsp112_42 sp112_42 sp113_42 11.551961
Rsn112_42 sn112_42 sn113_42 11.551961
Rsp112_43 sp112_43 sp113_43 11.551961
Rsn112_43 sn112_43 sn113_43 11.551961
Rsp112_44 sp112_44 sp113_44 11.551961
Rsn112_44 sn112_44 sn113_44 11.551961
Rsp112_45 sp112_45 sp113_45 11.551961
Rsn112_45 sn112_45 sn113_45 11.551961
Rsp112_46 sp112_46 sp113_46 11.551961
Rsn112_46 sn112_46 sn113_46 11.551961
Rsp112_47 sp112_47 sp113_47 11.551961
Rsn112_47 sn112_47 sn113_47 11.551961
Rsp112_48 sp112_48 sp113_48 11.551961
Rsn112_48 sn112_48 sn113_48 11.551961
Rsp112_49 sp112_49 sp113_49 11.551961
Rsn112_49 sn112_49 sn113_49 11.551961
Rsp112_50 sp112_50 sp113_50 11.551961
Rsn112_50 sn112_50 sn113_50 11.551961
Rsp112_51 sp112_51 sp113_51 11.551961
Rsn112_51 sn112_51 sn113_51 11.551961
Rsp112_52 sp112_52 sp113_52 11.551961
Rsn112_52 sn112_52 sn113_52 11.551961
Rsp112_53 sp112_53 sp113_53 11.551961
Rsn112_53 sn112_53 sn113_53 11.551961
Rsp112_54 sp112_54 sp113_54 11.551961
Rsn112_54 sn112_54 sn113_54 11.551961
Rsp112_55 sp112_55 sp113_55 11.551961
Rsn112_55 sn112_55 sn113_55 11.551961
Rsp112_56 sp112_56 sp113_56 11.551961
Rsn112_56 sn112_56 sn113_56 11.551961
Rsp112_57 sp112_57 sp113_57 11.551961
Rsn112_57 sn112_57 sn113_57 11.551961
Rsp112_58 sp112_58 sp113_58 11.551961
Rsn112_58 sn112_58 sn113_58 11.551961
Rsp112_59 sp112_59 sp113_59 11.551961
Rsn112_59 sn112_59 sn113_59 11.551961
Rsp112_60 sp112_60 sp113_60 11.551961
Rsn112_60 sn112_60 sn113_60 11.551961
Rsp112_61 sp112_61 sp113_61 11.551961
Rsn112_61 sn112_61 sn113_61 11.551961
Rsp112_62 sp112_62 sp113_62 11.551961
Rsn112_62 sn112_62 sn113_62 11.551961
Rsp112_63 sp112_63 sp113_63 11.551961
Rsn112_63 sn112_63 sn113_63 11.551961
Rsp112_64 sp112_64 sp113_64 11.551961
Rsn112_64 sn112_64 sn113_64 11.551961
Rsp112_65 sp112_65 sp113_65 11.551961
Rsn112_65 sn112_65 sn113_65 11.551961
Rsp112_66 sp112_66 sp113_66 11.551961
Rsn112_66 sn112_66 sn113_66 11.551961
Rsp112_67 sp112_67 sp113_67 11.551961
Rsn112_67 sn112_67 sn113_67 11.551961
Rsp112_68 sp112_68 sp113_68 11.551961
Rsn112_68 sn112_68 sn113_68 11.551961
Rsp112_69 sp112_69 sp113_69 11.551961
Rsn112_69 sn112_69 sn113_69 11.551961
Rsp112_70 sp112_70 sp113_70 11.551961
Rsn112_70 sn112_70 sn113_70 11.551961
Rsp112_71 sp112_71 sp113_71 11.551961
Rsn112_71 sn112_71 sn113_71 11.551961
Rsp112_72 sp112_72 sp113_72 11.551961
Rsn112_72 sn112_72 sn113_72 11.551961
Rsp112_73 sp112_73 sp113_73 11.551961
Rsn112_73 sn112_73 sn113_73 11.551961
Rsp112_74 sp112_74 sp113_74 11.551961
Rsn112_74 sn112_74 sn113_74 11.551961
Rsp112_75 sp112_75 sp113_75 11.551961
Rsn112_75 sn112_75 sn113_75 11.551961
Rsp112_76 sp112_76 sp113_76 11.551961
Rsn112_76 sn112_76 sn113_76 11.551961
Rsp112_77 sp112_77 sp113_77 11.551961
Rsn112_77 sn112_77 sn113_77 11.551961
Rsp112_78 sp112_78 sp113_78 11.551961
Rsn112_78 sn112_78 sn113_78 11.551961
Rsp112_79 sp112_79 sp113_79 11.551961
Rsn112_79 sn112_79 sn113_79 11.551961
Rsp112_80 sp112_80 sp113_80 11.551961
Rsn112_80 sn112_80 sn113_80 11.551961
Rsp112_81 sp112_81 sp113_81 11.551961
Rsn112_81 sn112_81 sn113_81 11.551961
Rsp112_82 sp112_82 sp113_82 11.551961
Rsn112_82 sn112_82 sn113_82 11.551961
Rsp112_83 sp112_83 sp113_83 11.551961
Rsn112_83 sn112_83 sn113_83 11.551961
Rsp112_84 sp112_84 sp113_84 11.551961
Rsn112_84 sn112_84 sn113_84 11.551961
Rsp113_1 sp113_1 sp114_1 11.551961
Rsn113_1 sn113_1 sn114_1 11.551961
Rsp113_2 sp113_2 sp114_2 11.551961
Rsn113_2 sn113_2 sn114_2 11.551961
Rsp113_3 sp113_3 sp114_3 11.551961
Rsn113_3 sn113_3 sn114_3 11.551961
Rsp113_4 sp113_4 sp114_4 11.551961
Rsn113_4 sn113_4 sn114_4 11.551961
Rsp113_5 sp113_5 sp114_5 11.551961
Rsn113_5 sn113_5 sn114_5 11.551961
Rsp113_6 sp113_6 sp114_6 11.551961
Rsn113_6 sn113_6 sn114_6 11.551961
Rsp113_7 sp113_7 sp114_7 11.551961
Rsn113_7 sn113_7 sn114_7 11.551961
Rsp113_8 sp113_8 sp114_8 11.551961
Rsn113_8 sn113_8 sn114_8 11.551961
Rsp113_9 sp113_9 sp114_9 11.551961
Rsn113_9 sn113_9 sn114_9 11.551961
Rsp113_10 sp113_10 sp114_10 11.551961
Rsn113_10 sn113_10 sn114_10 11.551961
Rsp113_11 sp113_11 sp114_11 11.551961
Rsn113_11 sn113_11 sn114_11 11.551961
Rsp113_12 sp113_12 sp114_12 11.551961
Rsn113_12 sn113_12 sn114_12 11.551961
Rsp113_13 sp113_13 sp114_13 11.551961
Rsn113_13 sn113_13 sn114_13 11.551961
Rsp113_14 sp113_14 sp114_14 11.551961
Rsn113_14 sn113_14 sn114_14 11.551961
Rsp113_15 sp113_15 sp114_15 11.551961
Rsn113_15 sn113_15 sn114_15 11.551961
Rsp113_16 sp113_16 sp114_16 11.551961
Rsn113_16 sn113_16 sn114_16 11.551961
Rsp113_17 sp113_17 sp114_17 11.551961
Rsn113_17 sn113_17 sn114_17 11.551961
Rsp113_18 sp113_18 sp114_18 11.551961
Rsn113_18 sn113_18 sn114_18 11.551961
Rsp113_19 sp113_19 sp114_19 11.551961
Rsn113_19 sn113_19 sn114_19 11.551961
Rsp113_20 sp113_20 sp114_20 11.551961
Rsn113_20 sn113_20 sn114_20 11.551961
Rsp113_21 sp113_21 sp114_21 11.551961
Rsn113_21 sn113_21 sn114_21 11.551961
Rsp113_22 sp113_22 sp114_22 11.551961
Rsn113_22 sn113_22 sn114_22 11.551961
Rsp113_23 sp113_23 sp114_23 11.551961
Rsn113_23 sn113_23 sn114_23 11.551961
Rsp113_24 sp113_24 sp114_24 11.551961
Rsn113_24 sn113_24 sn114_24 11.551961
Rsp113_25 sp113_25 sp114_25 11.551961
Rsn113_25 sn113_25 sn114_25 11.551961
Rsp113_26 sp113_26 sp114_26 11.551961
Rsn113_26 sn113_26 sn114_26 11.551961
Rsp113_27 sp113_27 sp114_27 11.551961
Rsn113_27 sn113_27 sn114_27 11.551961
Rsp113_28 sp113_28 sp114_28 11.551961
Rsn113_28 sn113_28 sn114_28 11.551961
Rsp113_29 sp113_29 sp114_29 11.551961
Rsn113_29 sn113_29 sn114_29 11.551961
Rsp113_30 sp113_30 sp114_30 11.551961
Rsn113_30 sn113_30 sn114_30 11.551961
Rsp113_31 sp113_31 sp114_31 11.551961
Rsn113_31 sn113_31 sn114_31 11.551961
Rsp113_32 sp113_32 sp114_32 11.551961
Rsn113_32 sn113_32 sn114_32 11.551961
Rsp113_33 sp113_33 sp114_33 11.551961
Rsn113_33 sn113_33 sn114_33 11.551961
Rsp113_34 sp113_34 sp114_34 11.551961
Rsn113_34 sn113_34 sn114_34 11.551961
Rsp113_35 sp113_35 sp114_35 11.551961
Rsn113_35 sn113_35 sn114_35 11.551961
Rsp113_36 sp113_36 sp114_36 11.551961
Rsn113_36 sn113_36 sn114_36 11.551961
Rsp113_37 sp113_37 sp114_37 11.551961
Rsn113_37 sn113_37 sn114_37 11.551961
Rsp113_38 sp113_38 sp114_38 11.551961
Rsn113_38 sn113_38 sn114_38 11.551961
Rsp113_39 sp113_39 sp114_39 11.551961
Rsn113_39 sn113_39 sn114_39 11.551961
Rsp113_40 sp113_40 sp114_40 11.551961
Rsn113_40 sn113_40 sn114_40 11.551961
Rsp113_41 sp113_41 sp114_41 11.551961
Rsn113_41 sn113_41 sn114_41 11.551961
Rsp113_42 sp113_42 sp114_42 11.551961
Rsn113_42 sn113_42 sn114_42 11.551961
Rsp113_43 sp113_43 sp114_43 11.551961
Rsn113_43 sn113_43 sn114_43 11.551961
Rsp113_44 sp113_44 sp114_44 11.551961
Rsn113_44 sn113_44 sn114_44 11.551961
Rsp113_45 sp113_45 sp114_45 11.551961
Rsn113_45 sn113_45 sn114_45 11.551961
Rsp113_46 sp113_46 sp114_46 11.551961
Rsn113_46 sn113_46 sn114_46 11.551961
Rsp113_47 sp113_47 sp114_47 11.551961
Rsn113_47 sn113_47 sn114_47 11.551961
Rsp113_48 sp113_48 sp114_48 11.551961
Rsn113_48 sn113_48 sn114_48 11.551961
Rsp113_49 sp113_49 sp114_49 11.551961
Rsn113_49 sn113_49 sn114_49 11.551961
Rsp113_50 sp113_50 sp114_50 11.551961
Rsn113_50 sn113_50 sn114_50 11.551961
Rsp113_51 sp113_51 sp114_51 11.551961
Rsn113_51 sn113_51 sn114_51 11.551961
Rsp113_52 sp113_52 sp114_52 11.551961
Rsn113_52 sn113_52 sn114_52 11.551961
Rsp113_53 sp113_53 sp114_53 11.551961
Rsn113_53 sn113_53 sn114_53 11.551961
Rsp113_54 sp113_54 sp114_54 11.551961
Rsn113_54 sn113_54 sn114_54 11.551961
Rsp113_55 sp113_55 sp114_55 11.551961
Rsn113_55 sn113_55 sn114_55 11.551961
Rsp113_56 sp113_56 sp114_56 11.551961
Rsn113_56 sn113_56 sn114_56 11.551961
Rsp113_57 sp113_57 sp114_57 11.551961
Rsn113_57 sn113_57 sn114_57 11.551961
Rsp113_58 sp113_58 sp114_58 11.551961
Rsn113_58 sn113_58 sn114_58 11.551961
Rsp113_59 sp113_59 sp114_59 11.551961
Rsn113_59 sn113_59 sn114_59 11.551961
Rsp113_60 sp113_60 sp114_60 11.551961
Rsn113_60 sn113_60 sn114_60 11.551961
Rsp113_61 sp113_61 sp114_61 11.551961
Rsn113_61 sn113_61 sn114_61 11.551961
Rsp113_62 sp113_62 sp114_62 11.551961
Rsn113_62 sn113_62 sn114_62 11.551961
Rsp113_63 sp113_63 sp114_63 11.551961
Rsn113_63 sn113_63 sn114_63 11.551961
Rsp113_64 sp113_64 sp114_64 11.551961
Rsn113_64 sn113_64 sn114_64 11.551961
Rsp113_65 sp113_65 sp114_65 11.551961
Rsn113_65 sn113_65 sn114_65 11.551961
Rsp113_66 sp113_66 sp114_66 11.551961
Rsn113_66 sn113_66 sn114_66 11.551961
Rsp113_67 sp113_67 sp114_67 11.551961
Rsn113_67 sn113_67 sn114_67 11.551961
Rsp113_68 sp113_68 sp114_68 11.551961
Rsn113_68 sn113_68 sn114_68 11.551961
Rsp113_69 sp113_69 sp114_69 11.551961
Rsn113_69 sn113_69 sn114_69 11.551961
Rsp113_70 sp113_70 sp114_70 11.551961
Rsn113_70 sn113_70 sn114_70 11.551961
Rsp113_71 sp113_71 sp114_71 11.551961
Rsn113_71 sn113_71 sn114_71 11.551961
Rsp113_72 sp113_72 sp114_72 11.551961
Rsn113_72 sn113_72 sn114_72 11.551961
Rsp113_73 sp113_73 sp114_73 11.551961
Rsn113_73 sn113_73 sn114_73 11.551961
Rsp113_74 sp113_74 sp114_74 11.551961
Rsn113_74 sn113_74 sn114_74 11.551961
Rsp113_75 sp113_75 sp114_75 11.551961
Rsn113_75 sn113_75 sn114_75 11.551961
Rsp113_76 sp113_76 sp114_76 11.551961
Rsn113_76 sn113_76 sn114_76 11.551961
Rsp113_77 sp113_77 sp114_77 11.551961
Rsn113_77 sn113_77 sn114_77 11.551961
Rsp113_78 sp113_78 sp114_78 11.551961
Rsn113_78 sn113_78 sn114_78 11.551961
Rsp113_79 sp113_79 sp114_79 11.551961
Rsn113_79 sn113_79 sn114_79 11.551961
Rsp113_80 sp113_80 sp114_80 11.551961
Rsn113_80 sn113_80 sn114_80 11.551961
Rsp113_81 sp113_81 sp114_81 11.551961
Rsn113_81 sn113_81 sn114_81 11.551961
Rsp113_82 sp113_82 sp114_82 11.551961
Rsn113_82 sn113_82 sn114_82 11.551961
Rsp113_83 sp113_83 sp114_83 11.551961
Rsn113_83 sn113_83 sn114_83 11.551961
Rsp113_84 sp113_84 sp114_84 11.551961
Rsn113_84 sn113_84 sn114_84 11.551961
Rsp114_1 sp114_1 sp115_1 11.551961
Rsn114_1 sn114_1 sn115_1 11.551961
Rsp114_2 sp114_2 sp115_2 11.551961
Rsn114_2 sn114_2 sn115_2 11.551961
Rsp114_3 sp114_3 sp115_3 11.551961
Rsn114_3 sn114_3 sn115_3 11.551961
Rsp114_4 sp114_4 sp115_4 11.551961
Rsn114_4 sn114_4 sn115_4 11.551961
Rsp114_5 sp114_5 sp115_5 11.551961
Rsn114_5 sn114_5 sn115_5 11.551961
Rsp114_6 sp114_6 sp115_6 11.551961
Rsn114_6 sn114_6 sn115_6 11.551961
Rsp114_7 sp114_7 sp115_7 11.551961
Rsn114_7 sn114_7 sn115_7 11.551961
Rsp114_8 sp114_8 sp115_8 11.551961
Rsn114_8 sn114_8 sn115_8 11.551961
Rsp114_9 sp114_9 sp115_9 11.551961
Rsn114_9 sn114_9 sn115_9 11.551961
Rsp114_10 sp114_10 sp115_10 11.551961
Rsn114_10 sn114_10 sn115_10 11.551961
Rsp114_11 sp114_11 sp115_11 11.551961
Rsn114_11 sn114_11 sn115_11 11.551961
Rsp114_12 sp114_12 sp115_12 11.551961
Rsn114_12 sn114_12 sn115_12 11.551961
Rsp114_13 sp114_13 sp115_13 11.551961
Rsn114_13 sn114_13 sn115_13 11.551961
Rsp114_14 sp114_14 sp115_14 11.551961
Rsn114_14 sn114_14 sn115_14 11.551961
Rsp114_15 sp114_15 sp115_15 11.551961
Rsn114_15 sn114_15 sn115_15 11.551961
Rsp114_16 sp114_16 sp115_16 11.551961
Rsn114_16 sn114_16 sn115_16 11.551961
Rsp114_17 sp114_17 sp115_17 11.551961
Rsn114_17 sn114_17 sn115_17 11.551961
Rsp114_18 sp114_18 sp115_18 11.551961
Rsn114_18 sn114_18 sn115_18 11.551961
Rsp114_19 sp114_19 sp115_19 11.551961
Rsn114_19 sn114_19 sn115_19 11.551961
Rsp114_20 sp114_20 sp115_20 11.551961
Rsn114_20 sn114_20 sn115_20 11.551961
Rsp114_21 sp114_21 sp115_21 11.551961
Rsn114_21 sn114_21 sn115_21 11.551961
Rsp114_22 sp114_22 sp115_22 11.551961
Rsn114_22 sn114_22 sn115_22 11.551961
Rsp114_23 sp114_23 sp115_23 11.551961
Rsn114_23 sn114_23 sn115_23 11.551961
Rsp114_24 sp114_24 sp115_24 11.551961
Rsn114_24 sn114_24 sn115_24 11.551961
Rsp114_25 sp114_25 sp115_25 11.551961
Rsn114_25 sn114_25 sn115_25 11.551961
Rsp114_26 sp114_26 sp115_26 11.551961
Rsn114_26 sn114_26 sn115_26 11.551961
Rsp114_27 sp114_27 sp115_27 11.551961
Rsn114_27 sn114_27 sn115_27 11.551961
Rsp114_28 sp114_28 sp115_28 11.551961
Rsn114_28 sn114_28 sn115_28 11.551961
Rsp114_29 sp114_29 sp115_29 11.551961
Rsn114_29 sn114_29 sn115_29 11.551961
Rsp114_30 sp114_30 sp115_30 11.551961
Rsn114_30 sn114_30 sn115_30 11.551961
Rsp114_31 sp114_31 sp115_31 11.551961
Rsn114_31 sn114_31 sn115_31 11.551961
Rsp114_32 sp114_32 sp115_32 11.551961
Rsn114_32 sn114_32 sn115_32 11.551961
Rsp114_33 sp114_33 sp115_33 11.551961
Rsn114_33 sn114_33 sn115_33 11.551961
Rsp114_34 sp114_34 sp115_34 11.551961
Rsn114_34 sn114_34 sn115_34 11.551961
Rsp114_35 sp114_35 sp115_35 11.551961
Rsn114_35 sn114_35 sn115_35 11.551961
Rsp114_36 sp114_36 sp115_36 11.551961
Rsn114_36 sn114_36 sn115_36 11.551961
Rsp114_37 sp114_37 sp115_37 11.551961
Rsn114_37 sn114_37 sn115_37 11.551961
Rsp114_38 sp114_38 sp115_38 11.551961
Rsn114_38 sn114_38 sn115_38 11.551961
Rsp114_39 sp114_39 sp115_39 11.551961
Rsn114_39 sn114_39 sn115_39 11.551961
Rsp114_40 sp114_40 sp115_40 11.551961
Rsn114_40 sn114_40 sn115_40 11.551961
Rsp114_41 sp114_41 sp115_41 11.551961
Rsn114_41 sn114_41 sn115_41 11.551961
Rsp114_42 sp114_42 sp115_42 11.551961
Rsn114_42 sn114_42 sn115_42 11.551961
Rsp114_43 sp114_43 sp115_43 11.551961
Rsn114_43 sn114_43 sn115_43 11.551961
Rsp114_44 sp114_44 sp115_44 11.551961
Rsn114_44 sn114_44 sn115_44 11.551961
Rsp114_45 sp114_45 sp115_45 11.551961
Rsn114_45 sn114_45 sn115_45 11.551961
Rsp114_46 sp114_46 sp115_46 11.551961
Rsn114_46 sn114_46 sn115_46 11.551961
Rsp114_47 sp114_47 sp115_47 11.551961
Rsn114_47 sn114_47 sn115_47 11.551961
Rsp114_48 sp114_48 sp115_48 11.551961
Rsn114_48 sn114_48 sn115_48 11.551961
Rsp114_49 sp114_49 sp115_49 11.551961
Rsn114_49 sn114_49 sn115_49 11.551961
Rsp114_50 sp114_50 sp115_50 11.551961
Rsn114_50 sn114_50 sn115_50 11.551961
Rsp114_51 sp114_51 sp115_51 11.551961
Rsn114_51 sn114_51 sn115_51 11.551961
Rsp114_52 sp114_52 sp115_52 11.551961
Rsn114_52 sn114_52 sn115_52 11.551961
Rsp114_53 sp114_53 sp115_53 11.551961
Rsn114_53 sn114_53 sn115_53 11.551961
Rsp114_54 sp114_54 sp115_54 11.551961
Rsn114_54 sn114_54 sn115_54 11.551961
Rsp114_55 sp114_55 sp115_55 11.551961
Rsn114_55 sn114_55 sn115_55 11.551961
Rsp114_56 sp114_56 sp115_56 11.551961
Rsn114_56 sn114_56 sn115_56 11.551961
Rsp114_57 sp114_57 sp115_57 11.551961
Rsn114_57 sn114_57 sn115_57 11.551961
Rsp114_58 sp114_58 sp115_58 11.551961
Rsn114_58 sn114_58 sn115_58 11.551961
Rsp114_59 sp114_59 sp115_59 11.551961
Rsn114_59 sn114_59 sn115_59 11.551961
Rsp114_60 sp114_60 sp115_60 11.551961
Rsn114_60 sn114_60 sn115_60 11.551961
Rsp114_61 sp114_61 sp115_61 11.551961
Rsn114_61 sn114_61 sn115_61 11.551961
Rsp114_62 sp114_62 sp115_62 11.551961
Rsn114_62 sn114_62 sn115_62 11.551961
Rsp114_63 sp114_63 sp115_63 11.551961
Rsn114_63 sn114_63 sn115_63 11.551961
Rsp114_64 sp114_64 sp115_64 11.551961
Rsn114_64 sn114_64 sn115_64 11.551961
Rsp114_65 sp114_65 sp115_65 11.551961
Rsn114_65 sn114_65 sn115_65 11.551961
Rsp114_66 sp114_66 sp115_66 11.551961
Rsn114_66 sn114_66 sn115_66 11.551961
Rsp114_67 sp114_67 sp115_67 11.551961
Rsn114_67 sn114_67 sn115_67 11.551961
Rsp114_68 sp114_68 sp115_68 11.551961
Rsn114_68 sn114_68 sn115_68 11.551961
Rsp114_69 sp114_69 sp115_69 11.551961
Rsn114_69 sn114_69 sn115_69 11.551961
Rsp114_70 sp114_70 sp115_70 11.551961
Rsn114_70 sn114_70 sn115_70 11.551961
Rsp114_71 sp114_71 sp115_71 11.551961
Rsn114_71 sn114_71 sn115_71 11.551961
Rsp114_72 sp114_72 sp115_72 11.551961
Rsn114_72 sn114_72 sn115_72 11.551961
Rsp114_73 sp114_73 sp115_73 11.551961
Rsn114_73 sn114_73 sn115_73 11.551961
Rsp114_74 sp114_74 sp115_74 11.551961
Rsn114_74 sn114_74 sn115_74 11.551961
Rsp114_75 sp114_75 sp115_75 11.551961
Rsn114_75 sn114_75 sn115_75 11.551961
Rsp114_76 sp114_76 sp115_76 11.551961
Rsn114_76 sn114_76 sn115_76 11.551961
Rsp114_77 sp114_77 sp115_77 11.551961
Rsn114_77 sn114_77 sn115_77 11.551961
Rsp114_78 sp114_78 sp115_78 11.551961
Rsn114_78 sn114_78 sn115_78 11.551961
Rsp114_79 sp114_79 sp115_79 11.551961
Rsn114_79 sn114_79 sn115_79 11.551961
Rsp114_80 sp114_80 sp115_80 11.551961
Rsn114_80 sn114_80 sn115_80 11.551961
Rsp114_81 sp114_81 sp115_81 11.551961
Rsn114_81 sn114_81 sn115_81 11.551961
Rsp114_82 sp114_82 sp115_82 11.551961
Rsn114_82 sn114_82 sn115_82 11.551961
Rsp114_83 sp114_83 sp115_83 11.551961
Rsn114_83 sn114_83 sn115_83 11.551961
Rsp114_84 sp114_84 sp115_84 11.551961
Rsn114_84 sn114_84 sn115_84 11.551961
Rsp115_1 sp115_1 sp116_1 11.551961
Rsn115_1 sn115_1 sn116_1 11.551961
Rsp115_2 sp115_2 sp116_2 11.551961
Rsn115_2 sn115_2 sn116_2 11.551961
Rsp115_3 sp115_3 sp116_3 11.551961
Rsn115_3 sn115_3 sn116_3 11.551961
Rsp115_4 sp115_4 sp116_4 11.551961
Rsn115_4 sn115_4 sn116_4 11.551961
Rsp115_5 sp115_5 sp116_5 11.551961
Rsn115_5 sn115_5 sn116_5 11.551961
Rsp115_6 sp115_6 sp116_6 11.551961
Rsn115_6 sn115_6 sn116_6 11.551961
Rsp115_7 sp115_7 sp116_7 11.551961
Rsn115_7 sn115_7 sn116_7 11.551961
Rsp115_8 sp115_8 sp116_8 11.551961
Rsn115_8 sn115_8 sn116_8 11.551961
Rsp115_9 sp115_9 sp116_9 11.551961
Rsn115_9 sn115_9 sn116_9 11.551961
Rsp115_10 sp115_10 sp116_10 11.551961
Rsn115_10 sn115_10 sn116_10 11.551961
Rsp115_11 sp115_11 sp116_11 11.551961
Rsn115_11 sn115_11 sn116_11 11.551961
Rsp115_12 sp115_12 sp116_12 11.551961
Rsn115_12 sn115_12 sn116_12 11.551961
Rsp115_13 sp115_13 sp116_13 11.551961
Rsn115_13 sn115_13 sn116_13 11.551961
Rsp115_14 sp115_14 sp116_14 11.551961
Rsn115_14 sn115_14 sn116_14 11.551961
Rsp115_15 sp115_15 sp116_15 11.551961
Rsn115_15 sn115_15 sn116_15 11.551961
Rsp115_16 sp115_16 sp116_16 11.551961
Rsn115_16 sn115_16 sn116_16 11.551961
Rsp115_17 sp115_17 sp116_17 11.551961
Rsn115_17 sn115_17 sn116_17 11.551961
Rsp115_18 sp115_18 sp116_18 11.551961
Rsn115_18 sn115_18 sn116_18 11.551961
Rsp115_19 sp115_19 sp116_19 11.551961
Rsn115_19 sn115_19 sn116_19 11.551961
Rsp115_20 sp115_20 sp116_20 11.551961
Rsn115_20 sn115_20 sn116_20 11.551961
Rsp115_21 sp115_21 sp116_21 11.551961
Rsn115_21 sn115_21 sn116_21 11.551961
Rsp115_22 sp115_22 sp116_22 11.551961
Rsn115_22 sn115_22 sn116_22 11.551961
Rsp115_23 sp115_23 sp116_23 11.551961
Rsn115_23 sn115_23 sn116_23 11.551961
Rsp115_24 sp115_24 sp116_24 11.551961
Rsn115_24 sn115_24 sn116_24 11.551961
Rsp115_25 sp115_25 sp116_25 11.551961
Rsn115_25 sn115_25 sn116_25 11.551961
Rsp115_26 sp115_26 sp116_26 11.551961
Rsn115_26 sn115_26 sn116_26 11.551961
Rsp115_27 sp115_27 sp116_27 11.551961
Rsn115_27 sn115_27 sn116_27 11.551961
Rsp115_28 sp115_28 sp116_28 11.551961
Rsn115_28 sn115_28 sn116_28 11.551961
Rsp115_29 sp115_29 sp116_29 11.551961
Rsn115_29 sn115_29 sn116_29 11.551961
Rsp115_30 sp115_30 sp116_30 11.551961
Rsn115_30 sn115_30 sn116_30 11.551961
Rsp115_31 sp115_31 sp116_31 11.551961
Rsn115_31 sn115_31 sn116_31 11.551961
Rsp115_32 sp115_32 sp116_32 11.551961
Rsn115_32 sn115_32 sn116_32 11.551961
Rsp115_33 sp115_33 sp116_33 11.551961
Rsn115_33 sn115_33 sn116_33 11.551961
Rsp115_34 sp115_34 sp116_34 11.551961
Rsn115_34 sn115_34 sn116_34 11.551961
Rsp115_35 sp115_35 sp116_35 11.551961
Rsn115_35 sn115_35 sn116_35 11.551961
Rsp115_36 sp115_36 sp116_36 11.551961
Rsn115_36 sn115_36 sn116_36 11.551961
Rsp115_37 sp115_37 sp116_37 11.551961
Rsn115_37 sn115_37 sn116_37 11.551961
Rsp115_38 sp115_38 sp116_38 11.551961
Rsn115_38 sn115_38 sn116_38 11.551961
Rsp115_39 sp115_39 sp116_39 11.551961
Rsn115_39 sn115_39 sn116_39 11.551961
Rsp115_40 sp115_40 sp116_40 11.551961
Rsn115_40 sn115_40 sn116_40 11.551961
Rsp115_41 sp115_41 sp116_41 11.551961
Rsn115_41 sn115_41 sn116_41 11.551961
Rsp115_42 sp115_42 sp116_42 11.551961
Rsn115_42 sn115_42 sn116_42 11.551961
Rsp115_43 sp115_43 sp116_43 11.551961
Rsn115_43 sn115_43 sn116_43 11.551961
Rsp115_44 sp115_44 sp116_44 11.551961
Rsn115_44 sn115_44 sn116_44 11.551961
Rsp115_45 sp115_45 sp116_45 11.551961
Rsn115_45 sn115_45 sn116_45 11.551961
Rsp115_46 sp115_46 sp116_46 11.551961
Rsn115_46 sn115_46 sn116_46 11.551961
Rsp115_47 sp115_47 sp116_47 11.551961
Rsn115_47 sn115_47 sn116_47 11.551961
Rsp115_48 sp115_48 sp116_48 11.551961
Rsn115_48 sn115_48 sn116_48 11.551961
Rsp115_49 sp115_49 sp116_49 11.551961
Rsn115_49 sn115_49 sn116_49 11.551961
Rsp115_50 sp115_50 sp116_50 11.551961
Rsn115_50 sn115_50 sn116_50 11.551961
Rsp115_51 sp115_51 sp116_51 11.551961
Rsn115_51 sn115_51 sn116_51 11.551961
Rsp115_52 sp115_52 sp116_52 11.551961
Rsn115_52 sn115_52 sn116_52 11.551961
Rsp115_53 sp115_53 sp116_53 11.551961
Rsn115_53 sn115_53 sn116_53 11.551961
Rsp115_54 sp115_54 sp116_54 11.551961
Rsn115_54 sn115_54 sn116_54 11.551961
Rsp115_55 sp115_55 sp116_55 11.551961
Rsn115_55 sn115_55 sn116_55 11.551961
Rsp115_56 sp115_56 sp116_56 11.551961
Rsn115_56 sn115_56 sn116_56 11.551961
Rsp115_57 sp115_57 sp116_57 11.551961
Rsn115_57 sn115_57 sn116_57 11.551961
Rsp115_58 sp115_58 sp116_58 11.551961
Rsn115_58 sn115_58 sn116_58 11.551961
Rsp115_59 sp115_59 sp116_59 11.551961
Rsn115_59 sn115_59 sn116_59 11.551961
Rsp115_60 sp115_60 sp116_60 11.551961
Rsn115_60 sn115_60 sn116_60 11.551961
Rsp115_61 sp115_61 sp116_61 11.551961
Rsn115_61 sn115_61 sn116_61 11.551961
Rsp115_62 sp115_62 sp116_62 11.551961
Rsn115_62 sn115_62 sn116_62 11.551961
Rsp115_63 sp115_63 sp116_63 11.551961
Rsn115_63 sn115_63 sn116_63 11.551961
Rsp115_64 sp115_64 sp116_64 11.551961
Rsn115_64 sn115_64 sn116_64 11.551961
Rsp115_65 sp115_65 sp116_65 11.551961
Rsn115_65 sn115_65 sn116_65 11.551961
Rsp115_66 sp115_66 sp116_66 11.551961
Rsn115_66 sn115_66 sn116_66 11.551961
Rsp115_67 sp115_67 sp116_67 11.551961
Rsn115_67 sn115_67 sn116_67 11.551961
Rsp115_68 sp115_68 sp116_68 11.551961
Rsn115_68 sn115_68 sn116_68 11.551961
Rsp115_69 sp115_69 sp116_69 11.551961
Rsn115_69 sn115_69 sn116_69 11.551961
Rsp115_70 sp115_70 sp116_70 11.551961
Rsn115_70 sn115_70 sn116_70 11.551961
Rsp115_71 sp115_71 sp116_71 11.551961
Rsn115_71 sn115_71 sn116_71 11.551961
Rsp115_72 sp115_72 sp116_72 11.551961
Rsn115_72 sn115_72 sn116_72 11.551961
Rsp115_73 sp115_73 sp116_73 11.551961
Rsn115_73 sn115_73 sn116_73 11.551961
Rsp115_74 sp115_74 sp116_74 11.551961
Rsn115_74 sn115_74 sn116_74 11.551961
Rsp115_75 sp115_75 sp116_75 11.551961
Rsn115_75 sn115_75 sn116_75 11.551961
Rsp115_76 sp115_76 sp116_76 11.551961
Rsn115_76 sn115_76 sn116_76 11.551961
Rsp115_77 sp115_77 sp116_77 11.551961
Rsn115_77 sn115_77 sn116_77 11.551961
Rsp115_78 sp115_78 sp116_78 11.551961
Rsn115_78 sn115_78 sn116_78 11.551961
Rsp115_79 sp115_79 sp116_79 11.551961
Rsn115_79 sn115_79 sn116_79 11.551961
Rsp115_80 sp115_80 sp116_80 11.551961
Rsn115_80 sn115_80 sn116_80 11.551961
Rsp115_81 sp115_81 sp116_81 11.551961
Rsn115_81 sn115_81 sn116_81 11.551961
Rsp115_82 sp115_82 sp116_82 11.551961
Rsn115_82 sn115_82 sn116_82 11.551961
Rsp115_83 sp115_83 sp116_83 11.551961
Rsn115_83 sn115_83 sn116_83 11.551961
Rsp115_84 sp115_84 sp116_84 11.551961
Rsn115_84 sn115_84 sn116_84 11.551961
Rsp116_1 sp116_1 sp117_1 11.551961
Rsn116_1 sn116_1 sn117_1 11.551961
Rsp116_2 sp116_2 sp117_2 11.551961
Rsn116_2 sn116_2 sn117_2 11.551961
Rsp116_3 sp116_3 sp117_3 11.551961
Rsn116_3 sn116_3 sn117_3 11.551961
Rsp116_4 sp116_4 sp117_4 11.551961
Rsn116_4 sn116_4 sn117_4 11.551961
Rsp116_5 sp116_5 sp117_5 11.551961
Rsn116_5 sn116_5 sn117_5 11.551961
Rsp116_6 sp116_6 sp117_6 11.551961
Rsn116_6 sn116_6 sn117_6 11.551961
Rsp116_7 sp116_7 sp117_7 11.551961
Rsn116_7 sn116_7 sn117_7 11.551961
Rsp116_8 sp116_8 sp117_8 11.551961
Rsn116_8 sn116_8 sn117_8 11.551961
Rsp116_9 sp116_9 sp117_9 11.551961
Rsn116_9 sn116_9 sn117_9 11.551961
Rsp116_10 sp116_10 sp117_10 11.551961
Rsn116_10 sn116_10 sn117_10 11.551961
Rsp116_11 sp116_11 sp117_11 11.551961
Rsn116_11 sn116_11 sn117_11 11.551961
Rsp116_12 sp116_12 sp117_12 11.551961
Rsn116_12 sn116_12 sn117_12 11.551961
Rsp116_13 sp116_13 sp117_13 11.551961
Rsn116_13 sn116_13 sn117_13 11.551961
Rsp116_14 sp116_14 sp117_14 11.551961
Rsn116_14 sn116_14 sn117_14 11.551961
Rsp116_15 sp116_15 sp117_15 11.551961
Rsn116_15 sn116_15 sn117_15 11.551961
Rsp116_16 sp116_16 sp117_16 11.551961
Rsn116_16 sn116_16 sn117_16 11.551961
Rsp116_17 sp116_17 sp117_17 11.551961
Rsn116_17 sn116_17 sn117_17 11.551961
Rsp116_18 sp116_18 sp117_18 11.551961
Rsn116_18 sn116_18 sn117_18 11.551961
Rsp116_19 sp116_19 sp117_19 11.551961
Rsn116_19 sn116_19 sn117_19 11.551961
Rsp116_20 sp116_20 sp117_20 11.551961
Rsn116_20 sn116_20 sn117_20 11.551961
Rsp116_21 sp116_21 sp117_21 11.551961
Rsn116_21 sn116_21 sn117_21 11.551961
Rsp116_22 sp116_22 sp117_22 11.551961
Rsn116_22 sn116_22 sn117_22 11.551961
Rsp116_23 sp116_23 sp117_23 11.551961
Rsn116_23 sn116_23 sn117_23 11.551961
Rsp116_24 sp116_24 sp117_24 11.551961
Rsn116_24 sn116_24 sn117_24 11.551961
Rsp116_25 sp116_25 sp117_25 11.551961
Rsn116_25 sn116_25 sn117_25 11.551961
Rsp116_26 sp116_26 sp117_26 11.551961
Rsn116_26 sn116_26 sn117_26 11.551961
Rsp116_27 sp116_27 sp117_27 11.551961
Rsn116_27 sn116_27 sn117_27 11.551961
Rsp116_28 sp116_28 sp117_28 11.551961
Rsn116_28 sn116_28 sn117_28 11.551961
Rsp116_29 sp116_29 sp117_29 11.551961
Rsn116_29 sn116_29 sn117_29 11.551961
Rsp116_30 sp116_30 sp117_30 11.551961
Rsn116_30 sn116_30 sn117_30 11.551961
Rsp116_31 sp116_31 sp117_31 11.551961
Rsn116_31 sn116_31 sn117_31 11.551961
Rsp116_32 sp116_32 sp117_32 11.551961
Rsn116_32 sn116_32 sn117_32 11.551961
Rsp116_33 sp116_33 sp117_33 11.551961
Rsn116_33 sn116_33 sn117_33 11.551961
Rsp116_34 sp116_34 sp117_34 11.551961
Rsn116_34 sn116_34 sn117_34 11.551961
Rsp116_35 sp116_35 sp117_35 11.551961
Rsn116_35 sn116_35 sn117_35 11.551961
Rsp116_36 sp116_36 sp117_36 11.551961
Rsn116_36 sn116_36 sn117_36 11.551961
Rsp116_37 sp116_37 sp117_37 11.551961
Rsn116_37 sn116_37 sn117_37 11.551961
Rsp116_38 sp116_38 sp117_38 11.551961
Rsn116_38 sn116_38 sn117_38 11.551961
Rsp116_39 sp116_39 sp117_39 11.551961
Rsn116_39 sn116_39 sn117_39 11.551961
Rsp116_40 sp116_40 sp117_40 11.551961
Rsn116_40 sn116_40 sn117_40 11.551961
Rsp116_41 sp116_41 sp117_41 11.551961
Rsn116_41 sn116_41 sn117_41 11.551961
Rsp116_42 sp116_42 sp117_42 11.551961
Rsn116_42 sn116_42 sn117_42 11.551961
Rsp116_43 sp116_43 sp117_43 11.551961
Rsn116_43 sn116_43 sn117_43 11.551961
Rsp116_44 sp116_44 sp117_44 11.551961
Rsn116_44 sn116_44 sn117_44 11.551961
Rsp116_45 sp116_45 sp117_45 11.551961
Rsn116_45 sn116_45 sn117_45 11.551961
Rsp116_46 sp116_46 sp117_46 11.551961
Rsn116_46 sn116_46 sn117_46 11.551961
Rsp116_47 sp116_47 sp117_47 11.551961
Rsn116_47 sn116_47 sn117_47 11.551961
Rsp116_48 sp116_48 sp117_48 11.551961
Rsn116_48 sn116_48 sn117_48 11.551961
Rsp116_49 sp116_49 sp117_49 11.551961
Rsn116_49 sn116_49 sn117_49 11.551961
Rsp116_50 sp116_50 sp117_50 11.551961
Rsn116_50 sn116_50 sn117_50 11.551961
Rsp116_51 sp116_51 sp117_51 11.551961
Rsn116_51 sn116_51 sn117_51 11.551961
Rsp116_52 sp116_52 sp117_52 11.551961
Rsn116_52 sn116_52 sn117_52 11.551961
Rsp116_53 sp116_53 sp117_53 11.551961
Rsn116_53 sn116_53 sn117_53 11.551961
Rsp116_54 sp116_54 sp117_54 11.551961
Rsn116_54 sn116_54 sn117_54 11.551961
Rsp116_55 sp116_55 sp117_55 11.551961
Rsn116_55 sn116_55 sn117_55 11.551961
Rsp116_56 sp116_56 sp117_56 11.551961
Rsn116_56 sn116_56 sn117_56 11.551961
Rsp116_57 sp116_57 sp117_57 11.551961
Rsn116_57 sn116_57 sn117_57 11.551961
Rsp116_58 sp116_58 sp117_58 11.551961
Rsn116_58 sn116_58 sn117_58 11.551961
Rsp116_59 sp116_59 sp117_59 11.551961
Rsn116_59 sn116_59 sn117_59 11.551961
Rsp116_60 sp116_60 sp117_60 11.551961
Rsn116_60 sn116_60 sn117_60 11.551961
Rsp116_61 sp116_61 sp117_61 11.551961
Rsn116_61 sn116_61 sn117_61 11.551961
Rsp116_62 sp116_62 sp117_62 11.551961
Rsn116_62 sn116_62 sn117_62 11.551961
Rsp116_63 sp116_63 sp117_63 11.551961
Rsn116_63 sn116_63 sn117_63 11.551961
Rsp116_64 sp116_64 sp117_64 11.551961
Rsn116_64 sn116_64 sn117_64 11.551961
Rsp116_65 sp116_65 sp117_65 11.551961
Rsn116_65 sn116_65 sn117_65 11.551961
Rsp116_66 sp116_66 sp117_66 11.551961
Rsn116_66 sn116_66 sn117_66 11.551961
Rsp116_67 sp116_67 sp117_67 11.551961
Rsn116_67 sn116_67 sn117_67 11.551961
Rsp116_68 sp116_68 sp117_68 11.551961
Rsn116_68 sn116_68 sn117_68 11.551961
Rsp116_69 sp116_69 sp117_69 11.551961
Rsn116_69 sn116_69 sn117_69 11.551961
Rsp116_70 sp116_70 sp117_70 11.551961
Rsn116_70 sn116_70 sn117_70 11.551961
Rsp116_71 sp116_71 sp117_71 11.551961
Rsn116_71 sn116_71 sn117_71 11.551961
Rsp116_72 sp116_72 sp117_72 11.551961
Rsn116_72 sn116_72 sn117_72 11.551961
Rsp116_73 sp116_73 sp117_73 11.551961
Rsn116_73 sn116_73 sn117_73 11.551961
Rsp116_74 sp116_74 sp117_74 11.551961
Rsn116_74 sn116_74 sn117_74 11.551961
Rsp116_75 sp116_75 sp117_75 11.551961
Rsn116_75 sn116_75 sn117_75 11.551961
Rsp116_76 sp116_76 sp117_76 11.551961
Rsn116_76 sn116_76 sn117_76 11.551961
Rsp116_77 sp116_77 sp117_77 11.551961
Rsn116_77 sn116_77 sn117_77 11.551961
Rsp116_78 sp116_78 sp117_78 11.551961
Rsn116_78 sn116_78 sn117_78 11.551961
Rsp116_79 sp116_79 sp117_79 11.551961
Rsn116_79 sn116_79 sn117_79 11.551961
Rsp116_80 sp116_80 sp117_80 11.551961
Rsn116_80 sn116_80 sn117_80 11.551961
Rsp116_81 sp116_81 sp117_81 11.551961
Rsn116_81 sn116_81 sn117_81 11.551961
Rsp116_82 sp116_82 sp117_82 11.551961
Rsn116_82 sn116_82 sn117_82 11.551961
Rsp116_83 sp116_83 sp117_83 11.551961
Rsn116_83 sn116_83 sn117_83 11.551961
Rsp116_84 sp116_84 sp117_84 11.551961
Rsn116_84 sn116_84 sn117_84 11.551961
Rsp117_1 sp117_1 sp118_1 11.551961
Rsn117_1 sn117_1 sn118_1 11.551961
Rsp117_2 sp117_2 sp118_2 11.551961
Rsn117_2 sn117_2 sn118_2 11.551961
Rsp117_3 sp117_3 sp118_3 11.551961
Rsn117_3 sn117_3 sn118_3 11.551961
Rsp117_4 sp117_4 sp118_4 11.551961
Rsn117_4 sn117_4 sn118_4 11.551961
Rsp117_5 sp117_5 sp118_5 11.551961
Rsn117_5 sn117_5 sn118_5 11.551961
Rsp117_6 sp117_6 sp118_6 11.551961
Rsn117_6 sn117_6 sn118_6 11.551961
Rsp117_7 sp117_7 sp118_7 11.551961
Rsn117_7 sn117_7 sn118_7 11.551961
Rsp117_8 sp117_8 sp118_8 11.551961
Rsn117_8 sn117_8 sn118_8 11.551961
Rsp117_9 sp117_9 sp118_9 11.551961
Rsn117_9 sn117_9 sn118_9 11.551961
Rsp117_10 sp117_10 sp118_10 11.551961
Rsn117_10 sn117_10 sn118_10 11.551961
Rsp117_11 sp117_11 sp118_11 11.551961
Rsn117_11 sn117_11 sn118_11 11.551961
Rsp117_12 sp117_12 sp118_12 11.551961
Rsn117_12 sn117_12 sn118_12 11.551961
Rsp117_13 sp117_13 sp118_13 11.551961
Rsn117_13 sn117_13 sn118_13 11.551961
Rsp117_14 sp117_14 sp118_14 11.551961
Rsn117_14 sn117_14 sn118_14 11.551961
Rsp117_15 sp117_15 sp118_15 11.551961
Rsn117_15 sn117_15 sn118_15 11.551961
Rsp117_16 sp117_16 sp118_16 11.551961
Rsn117_16 sn117_16 sn118_16 11.551961
Rsp117_17 sp117_17 sp118_17 11.551961
Rsn117_17 sn117_17 sn118_17 11.551961
Rsp117_18 sp117_18 sp118_18 11.551961
Rsn117_18 sn117_18 sn118_18 11.551961
Rsp117_19 sp117_19 sp118_19 11.551961
Rsn117_19 sn117_19 sn118_19 11.551961
Rsp117_20 sp117_20 sp118_20 11.551961
Rsn117_20 sn117_20 sn118_20 11.551961
Rsp117_21 sp117_21 sp118_21 11.551961
Rsn117_21 sn117_21 sn118_21 11.551961
Rsp117_22 sp117_22 sp118_22 11.551961
Rsn117_22 sn117_22 sn118_22 11.551961
Rsp117_23 sp117_23 sp118_23 11.551961
Rsn117_23 sn117_23 sn118_23 11.551961
Rsp117_24 sp117_24 sp118_24 11.551961
Rsn117_24 sn117_24 sn118_24 11.551961
Rsp117_25 sp117_25 sp118_25 11.551961
Rsn117_25 sn117_25 sn118_25 11.551961
Rsp117_26 sp117_26 sp118_26 11.551961
Rsn117_26 sn117_26 sn118_26 11.551961
Rsp117_27 sp117_27 sp118_27 11.551961
Rsn117_27 sn117_27 sn118_27 11.551961
Rsp117_28 sp117_28 sp118_28 11.551961
Rsn117_28 sn117_28 sn118_28 11.551961
Rsp117_29 sp117_29 sp118_29 11.551961
Rsn117_29 sn117_29 sn118_29 11.551961
Rsp117_30 sp117_30 sp118_30 11.551961
Rsn117_30 sn117_30 sn118_30 11.551961
Rsp117_31 sp117_31 sp118_31 11.551961
Rsn117_31 sn117_31 sn118_31 11.551961
Rsp117_32 sp117_32 sp118_32 11.551961
Rsn117_32 sn117_32 sn118_32 11.551961
Rsp117_33 sp117_33 sp118_33 11.551961
Rsn117_33 sn117_33 sn118_33 11.551961
Rsp117_34 sp117_34 sp118_34 11.551961
Rsn117_34 sn117_34 sn118_34 11.551961
Rsp117_35 sp117_35 sp118_35 11.551961
Rsn117_35 sn117_35 sn118_35 11.551961
Rsp117_36 sp117_36 sp118_36 11.551961
Rsn117_36 sn117_36 sn118_36 11.551961
Rsp117_37 sp117_37 sp118_37 11.551961
Rsn117_37 sn117_37 sn118_37 11.551961
Rsp117_38 sp117_38 sp118_38 11.551961
Rsn117_38 sn117_38 sn118_38 11.551961
Rsp117_39 sp117_39 sp118_39 11.551961
Rsn117_39 sn117_39 sn118_39 11.551961
Rsp117_40 sp117_40 sp118_40 11.551961
Rsn117_40 sn117_40 sn118_40 11.551961
Rsp117_41 sp117_41 sp118_41 11.551961
Rsn117_41 sn117_41 sn118_41 11.551961
Rsp117_42 sp117_42 sp118_42 11.551961
Rsn117_42 sn117_42 sn118_42 11.551961
Rsp117_43 sp117_43 sp118_43 11.551961
Rsn117_43 sn117_43 sn118_43 11.551961
Rsp117_44 sp117_44 sp118_44 11.551961
Rsn117_44 sn117_44 sn118_44 11.551961
Rsp117_45 sp117_45 sp118_45 11.551961
Rsn117_45 sn117_45 sn118_45 11.551961
Rsp117_46 sp117_46 sp118_46 11.551961
Rsn117_46 sn117_46 sn118_46 11.551961
Rsp117_47 sp117_47 sp118_47 11.551961
Rsn117_47 sn117_47 sn118_47 11.551961
Rsp117_48 sp117_48 sp118_48 11.551961
Rsn117_48 sn117_48 sn118_48 11.551961
Rsp117_49 sp117_49 sp118_49 11.551961
Rsn117_49 sn117_49 sn118_49 11.551961
Rsp117_50 sp117_50 sp118_50 11.551961
Rsn117_50 sn117_50 sn118_50 11.551961
Rsp117_51 sp117_51 sp118_51 11.551961
Rsn117_51 sn117_51 sn118_51 11.551961
Rsp117_52 sp117_52 sp118_52 11.551961
Rsn117_52 sn117_52 sn118_52 11.551961
Rsp117_53 sp117_53 sp118_53 11.551961
Rsn117_53 sn117_53 sn118_53 11.551961
Rsp117_54 sp117_54 sp118_54 11.551961
Rsn117_54 sn117_54 sn118_54 11.551961
Rsp117_55 sp117_55 sp118_55 11.551961
Rsn117_55 sn117_55 sn118_55 11.551961
Rsp117_56 sp117_56 sp118_56 11.551961
Rsn117_56 sn117_56 sn118_56 11.551961
Rsp117_57 sp117_57 sp118_57 11.551961
Rsn117_57 sn117_57 sn118_57 11.551961
Rsp117_58 sp117_58 sp118_58 11.551961
Rsn117_58 sn117_58 sn118_58 11.551961
Rsp117_59 sp117_59 sp118_59 11.551961
Rsn117_59 sn117_59 sn118_59 11.551961
Rsp117_60 sp117_60 sp118_60 11.551961
Rsn117_60 sn117_60 sn118_60 11.551961
Rsp117_61 sp117_61 sp118_61 11.551961
Rsn117_61 sn117_61 sn118_61 11.551961
Rsp117_62 sp117_62 sp118_62 11.551961
Rsn117_62 sn117_62 sn118_62 11.551961
Rsp117_63 sp117_63 sp118_63 11.551961
Rsn117_63 sn117_63 sn118_63 11.551961
Rsp117_64 sp117_64 sp118_64 11.551961
Rsn117_64 sn117_64 sn118_64 11.551961
Rsp117_65 sp117_65 sp118_65 11.551961
Rsn117_65 sn117_65 sn118_65 11.551961
Rsp117_66 sp117_66 sp118_66 11.551961
Rsn117_66 sn117_66 sn118_66 11.551961
Rsp117_67 sp117_67 sp118_67 11.551961
Rsn117_67 sn117_67 sn118_67 11.551961
Rsp117_68 sp117_68 sp118_68 11.551961
Rsn117_68 sn117_68 sn118_68 11.551961
Rsp117_69 sp117_69 sp118_69 11.551961
Rsn117_69 sn117_69 sn118_69 11.551961
Rsp117_70 sp117_70 sp118_70 11.551961
Rsn117_70 sn117_70 sn118_70 11.551961
Rsp117_71 sp117_71 sp118_71 11.551961
Rsn117_71 sn117_71 sn118_71 11.551961
Rsp117_72 sp117_72 sp118_72 11.551961
Rsn117_72 sn117_72 sn118_72 11.551961
Rsp117_73 sp117_73 sp118_73 11.551961
Rsn117_73 sn117_73 sn118_73 11.551961
Rsp117_74 sp117_74 sp118_74 11.551961
Rsn117_74 sn117_74 sn118_74 11.551961
Rsp117_75 sp117_75 sp118_75 11.551961
Rsn117_75 sn117_75 sn118_75 11.551961
Rsp117_76 sp117_76 sp118_76 11.551961
Rsn117_76 sn117_76 sn118_76 11.551961
Rsp117_77 sp117_77 sp118_77 11.551961
Rsn117_77 sn117_77 sn118_77 11.551961
Rsp117_78 sp117_78 sp118_78 11.551961
Rsn117_78 sn117_78 sn118_78 11.551961
Rsp117_79 sp117_79 sp118_79 11.551961
Rsn117_79 sn117_79 sn118_79 11.551961
Rsp117_80 sp117_80 sp118_80 11.551961
Rsn117_80 sn117_80 sn118_80 11.551961
Rsp117_81 sp117_81 sp118_81 11.551961
Rsn117_81 sn117_81 sn118_81 11.551961
Rsp117_82 sp117_82 sp118_82 11.551961
Rsn117_82 sn117_82 sn118_82 11.551961
Rsp117_83 sp117_83 sp118_83 11.551961
Rsn117_83 sn117_83 sn118_83 11.551961
Rsp117_84 sp117_84 sp118_84 11.551961
Rsn117_84 sn117_84 sn118_84 11.551961
Rsp118_1 sp118_1 sp119_1 11.551961
Rsn118_1 sn118_1 sn119_1 11.551961
Rsp118_2 sp118_2 sp119_2 11.551961
Rsn118_2 sn118_2 sn119_2 11.551961
Rsp118_3 sp118_3 sp119_3 11.551961
Rsn118_3 sn118_3 sn119_3 11.551961
Rsp118_4 sp118_4 sp119_4 11.551961
Rsn118_4 sn118_4 sn119_4 11.551961
Rsp118_5 sp118_5 sp119_5 11.551961
Rsn118_5 sn118_5 sn119_5 11.551961
Rsp118_6 sp118_6 sp119_6 11.551961
Rsn118_6 sn118_6 sn119_6 11.551961
Rsp118_7 sp118_7 sp119_7 11.551961
Rsn118_7 sn118_7 sn119_7 11.551961
Rsp118_8 sp118_8 sp119_8 11.551961
Rsn118_8 sn118_8 sn119_8 11.551961
Rsp118_9 sp118_9 sp119_9 11.551961
Rsn118_9 sn118_9 sn119_9 11.551961
Rsp118_10 sp118_10 sp119_10 11.551961
Rsn118_10 sn118_10 sn119_10 11.551961
Rsp118_11 sp118_11 sp119_11 11.551961
Rsn118_11 sn118_11 sn119_11 11.551961
Rsp118_12 sp118_12 sp119_12 11.551961
Rsn118_12 sn118_12 sn119_12 11.551961
Rsp118_13 sp118_13 sp119_13 11.551961
Rsn118_13 sn118_13 sn119_13 11.551961
Rsp118_14 sp118_14 sp119_14 11.551961
Rsn118_14 sn118_14 sn119_14 11.551961
Rsp118_15 sp118_15 sp119_15 11.551961
Rsn118_15 sn118_15 sn119_15 11.551961
Rsp118_16 sp118_16 sp119_16 11.551961
Rsn118_16 sn118_16 sn119_16 11.551961
Rsp118_17 sp118_17 sp119_17 11.551961
Rsn118_17 sn118_17 sn119_17 11.551961
Rsp118_18 sp118_18 sp119_18 11.551961
Rsn118_18 sn118_18 sn119_18 11.551961
Rsp118_19 sp118_19 sp119_19 11.551961
Rsn118_19 sn118_19 sn119_19 11.551961
Rsp118_20 sp118_20 sp119_20 11.551961
Rsn118_20 sn118_20 sn119_20 11.551961
Rsp118_21 sp118_21 sp119_21 11.551961
Rsn118_21 sn118_21 sn119_21 11.551961
Rsp118_22 sp118_22 sp119_22 11.551961
Rsn118_22 sn118_22 sn119_22 11.551961
Rsp118_23 sp118_23 sp119_23 11.551961
Rsn118_23 sn118_23 sn119_23 11.551961
Rsp118_24 sp118_24 sp119_24 11.551961
Rsn118_24 sn118_24 sn119_24 11.551961
Rsp118_25 sp118_25 sp119_25 11.551961
Rsn118_25 sn118_25 sn119_25 11.551961
Rsp118_26 sp118_26 sp119_26 11.551961
Rsn118_26 sn118_26 sn119_26 11.551961
Rsp118_27 sp118_27 sp119_27 11.551961
Rsn118_27 sn118_27 sn119_27 11.551961
Rsp118_28 sp118_28 sp119_28 11.551961
Rsn118_28 sn118_28 sn119_28 11.551961
Rsp118_29 sp118_29 sp119_29 11.551961
Rsn118_29 sn118_29 sn119_29 11.551961
Rsp118_30 sp118_30 sp119_30 11.551961
Rsn118_30 sn118_30 sn119_30 11.551961
Rsp118_31 sp118_31 sp119_31 11.551961
Rsn118_31 sn118_31 sn119_31 11.551961
Rsp118_32 sp118_32 sp119_32 11.551961
Rsn118_32 sn118_32 sn119_32 11.551961
Rsp118_33 sp118_33 sp119_33 11.551961
Rsn118_33 sn118_33 sn119_33 11.551961
Rsp118_34 sp118_34 sp119_34 11.551961
Rsn118_34 sn118_34 sn119_34 11.551961
Rsp118_35 sp118_35 sp119_35 11.551961
Rsn118_35 sn118_35 sn119_35 11.551961
Rsp118_36 sp118_36 sp119_36 11.551961
Rsn118_36 sn118_36 sn119_36 11.551961
Rsp118_37 sp118_37 sp119_37 11.551961
Rsn118_37 sn118_37 sn119_37 11.551961
Rsp118_38 sp118_38 sp119_38 11.551961
Rsn118_38 sn118_38 sn119_38 11.551961
Rsp118_39 sp118_39 sp119_39 11.551961
Rsn118_39 sn118_39 sn119_39 11.551961
Rsp118_40 sp118_40 sp119_40 11.551961
Rsn118_40 sn118_40 sn119_40 11.551961
Rsp118_41 sp118_41 sp119_41 11.551961
Rsn118_41 sn118_41 sn119_41 11.551961
Rsp118_42 sp118_42 sp119_42 11.551961
Rsn118_42 sn118_42 sn119_42 11.551961
Rsp118_43 sp118_43 sp119_43 11.551961
Rsn118_43 sn118_43 sn119_43 11.551961
Rsp118_44 sp118_44 sp119_44 11.551961
Rsn118_44 sn118_44 sn119_44 11.551961
Rsp118_45 sp118_45 sp119_45 11.551961
Rsn118_45 sn118_45 sn119_45 11.551961
Rsp118_46 sp118_46 sp119_46 11.551961
Rsn118_46 sn118_46 sn119_46 11.551961
Rsp118_47 sp118_47 sp119_47 11.551961
Rsn118_47 sn118_47 sn119_47 11.551961
Rsp118_48 sp118_48 sp119_48 11.551961
Rsn118_48 sn118_48 sn119_48 11.551961
Rsp118_49 sp118_49 sp119_49 11.551961
Rsn118_49 sn118_49 sn119_49 11.551961
Rsp118_50 sp118_50 sp119_50 11.551961
Rsn118_50 sn118_50 sn119_50 11.551961
Rsp118_51 sp118_51 sp119_51 11.551961
Rsn118_51 sn118_51 sn119_51 11.551961
Rsp118_52 sp118_52 sp119_52 11.551961
Rsn118_52 sn118_52 sn119_52 11.551961
Rsp118_53 sp118_53 sp119_53 11.551961
Rsn118_53 sn118_53 sn119_53 11.551961
Rsp118_54 sp118_54 sp119_54 11.551961
Rsn118_54 sn118_54 sn119_54 11.551961
Rsp118_55 sp118_55 sp119_55 11.551961
Rsn118_55 sn118_55 sn119_55 11.551961
Rsp118_56 sp118_56 sp119_56 11.551961
Rsn118_56 sn118_56 sn119_56 11.551961
Rsp118_57 sp118_57 sp119_57 11.551961
Rsn118_57 sn118_57 sn119_57 11.551961
Rsp118_58 sp118_58 sp119_58 11.551961
Rsn118_58 sn118_58 sn119_58 11.551961
Rsp118_59 sp118_59 sp119_59 11.551961
Rsn118_59 sn118_59 sn119_59 11.551961
Rsp118_60 sp118_60 sp119_60 11.551961
Rsn118_60 sn118_60 sn119_60 11.551961
Rsp118_61 sp118_61 sp119_61 11.551961
Rsn118_61 sn118_61 sn119_61 11.551961
Rsp118_62 sp118_62 sp119_62 11.551961
Rsn118_62 sn118_62 sn119_62 11.551961
Rsp118_63 sp118_63 sp119_63 11.551961
Rsn118_63 sn118_63 sn119_63 11.551961
Rsp118_64 sp118_64 sp119_64 11.551961
Rsn118_64 sn118_64 sn119_64 11.551961
Rsp118_65 sp118_65 sp119_65 11.551961
Rsn118_65 sn118_65 sn119_65 11.551961
Rsp118_66 sp118_66 sp119_66 11.551961
Rsn118_66 sn118_66 sn119_66 11.551961
Rsp118_67 sp118_67 sp119_67 11.551961
Rsn118_67 sn118_67 sn119_67 11.551961
Rsp118_68 sp118_68 sp119_68 11.551961
Rsn118_68 sn118_68 sn119_68 11.551961
Rsp118_69 sp118_69 sp119_69 11.551961
Rsn118_69 sn118_69 sn119_69 11.551961
Rsp118_70 sp118_70 sp119_70 11.551961
Rsn118_70 sn118_70 sn119_70 11.551961
Rsp118_71 sp118_71 sp119_71 11.551961
Rsn118_71 sn118_71 sn119_71 11.551961
Rsp118_72 sp118_72 sp119_72 11.551961
Rsn118_72 sn118_72 sn119_72 11.551961
Rsp118_73 sp118_73 sp119_73 11.551961
Rsn118_73 sn118_73 sn119_73 11.551961
Rsp118_74 sp118_74 sp119_74 11.551961
Rsn118_74 sn118_74 sn119_74 11.551961
Rsp118_75 sp118_75 sp119_75 11.551961
Rsn118_75 sn118_75 sn119_75 11.551961
Rsp118_76 sp118_76 sp119_76 11.551961
Rsn118_76 sn118_76 sn119_76 11.551961
Rsp118_77 sp118_77 sp119_77 11.551961
Rsn118_77 sn118_77 sn119_77 11.551961
Rsp118_78 sp118_78 sp119_78 11.551961
Rsn118_78 sn118_78 sn119_78 11.551961
Rsp118_79 sp118_79 sp119_79 11.551961
Rsn118_79 sn118_79 sn119_79 11.551961
Rsp118_80 sp118_80 sp119_80 11.551961
Rsn118_80 sn118_80 sn119_80 11.551961
Rsp118_81 sp118_81 sp119_81 11.551961
Rsn118_81 sn118_81 sn119_81 11.551961
Rsp118_82 sp118_82 sp119_82 11.551961
Rsn118_82 sn118_82 sn119_82 11.551961
Rsp118_83 sp118_83 sp119_83 11.551961
Rsn118_83 sn118_83 sn119_83 11.551961
Rsp118_84 sp118_84 sp119_84 11.551961
Rsn118_84 sn118_84 sn119_84 11.551961
Rsp119_1 sp119_1 sp120_1 11.551961
Rsn119_1 sn119_1 sn120_1 11.551961
Rsp119_2 sp119_2 sp120_2 11.551961
Rsn119_2 sn119_2 sn120_2 11.551961
Rsp119_3 sp119_3 sp120_3 11.551961
Rsn119_3 sn119_3 sn120_3 11.551961
Rsp119_4 sp119_4 sp120_4 11.551961
Rsn119_4 sn119_4 sn120_4 11.551961
Rsp119_5 sp119_5 sp120_5 11.551961
Rsn119_5 sn119_5 sn120_5 11.551961
Rsp119_6 sp119_6 sp120_6 11.551961
Rsn119_6 sn119_6 sn120_6 11.551961
Rsp119_7 sp119_7 sp120_7 11.551961
Rsn119_7 sn119_7 sn120_7 11.551961
Rsp119_8 sp119_8 sp120_8 11.551961
Rsn119_8 sn119_8 sn120_8 11.551961
Rsp119_9 sp119_9 sp120_9 11.551961
Rsn119_9 sn119_9 sn120_9 11.551961
Rsp119_10 sp119_10 sp120_10 11.551961
Rsn119_10 sn119_10 sn120_10 11.551961
Rsp119_11 sp119_11 sp120_11 11.551961
Rsn119_11 sn119_11 sn120_11 11.551961
Rsp119_12 sp119_12 sp120_12 11.551961
Rsn119_12 sn119_12 sn120_12 11.551961
Rsp119_13 sp119_13 sp120_13 11.551961
Rsn119_13 sn119_13 sn120_13 11.551961
Rsp119_14 sp119_14 sp120_14 11.551961
Rsn119_14 sn119_14 sn120_14 11.551961
Rsp119_15 sp119_15 sp120_15 11.551961
Rsn119_15 sn119_15 sn120_15 11.551961
Rsp119_16 sp119_16 sp120_16 11.551961
Rsn119_16 sn119_16 sn120_16 11.551961
Rsp119_17 sp119_17 sp120_17 11.551961
Rsn119_17 sn119_17 sn120_17 11.551961
Rsp119_18 sp119_18 sp120_18 11.551961
Rsn119_18 sn119_18 sn120_18 11.551961
Rsp119_19 sp119_19 sp120_19 11.551961
Rsn119_19 sn119_19 sn120_19 11.551961
Rsp119_20 sp119_20 sp120_20 11.551961
Rsn119_20 sn119_20 sn120_20 11.551961
Rsp119_21 sp119_21 sp120_21 11.551961
Rsn119_21 sn119_21 sn120_21 11.551961
Rsp119_22 sp119_22 sp120_22 11.551961
Rsn119_22 sn119_22 sn120_22 11.551961
Rsp119_23 sp119_23 sp120_23 11.551961
Rsn119_23 sn119_23 sn120_23 11.551961
Rsp119_24 sp119_24 sp120_24 11.551961
Rsn119_24 sn119_24 sn120_24 11.551961
Rsp119_25 sp119_25 sp120_25 11.551961
Rsn119_25 sn119_25 sn120_25 11.551961
Rsp119_26 sp119_26 sp120_26 11.551961
Rsn119_26 sn119_26 sn120_26 11.551961
Rsp119_27 sp119_27 sp120_27 11.551961
Rsn119_27 sn119_27 sn120_27 11.551961
Rsp119_28 sp119_28 sp120_28 11.551961
Rsn119_28 sn119_28 sn120_28 11.551961
Rsp119_29 sp119_29 sp120_29 11.551961
Rsn119_29 sn119_29 sn120_29 11.551961
Rsp119_30 sp119_30 sp120_30 11.551961
Rsn119_30 sn119_30 sn120_30 11.551961
Rsp119_31 sp119_31 sp120_31 11.551961
Rsn119_31 sn119_31 sn120_31 11.551961
Rsp119_32 sp119_32 sp120_32 11.551961
Rsn119_32 sn119_32 sn120_32 11.551961
Rsp119_33 sp119_33 sp120_33 11.551961
Rsn119_33 sn119_33 sn120_33 11.551961
Rsp119_34 sp119_34 sp120_34 11.551961
Rsn119_34 sn119_34 sn120_34 11.551961
Rsp119_35 sp119_35 sp120_35 11.551961
Rsn119_35 sn119_35 sn120_35 11.551961
Rsp119_36 sp119_36 sp120_36 11.551961
Rsn119_36 sn119_36 sn120_36 11.551961
Rsp119_37 sp119_37 sp120_37 11.551961
Rsn119_37 sn119_37 sn120_37 11.551961
Rsp119_38 sp119_38 sp120_38 11.551961
Rsn119_38 sn119_38 sn120_38 11.551961
Rsp119_39 sp119_39 sp120_39 11.551961
Rsn119_39 sn119_39 sn120_39 11.551961
Rsp119_40 sp119_40 sp120_40 11.551961
Rsn119_40 sn119_40 sn120_40 11.551961
Rsp119_41 sp119_41 sp120_41 11.551961
Rsn119_41 sn119_41 sn120_41 11.551961
Rsp119_42 sp119_42 sp120_42 11.551961
Rsn119_42 sn119_42 sn120_42 11.551961
Rsp119_43 sp119_43 sp120_43 11.551961
Rsn119_43 sn119_43 sn120_43 11.551961
Rsp119_44 sp119_44 sp120_44 11.551961
Rsn119_44 sn119_44 sn120_44 11.551961
Rsp119_45 sp119_45 sp120_45 11.551961
Rsn119_45 sn119_45 sn120_45 11.551961
Rsp119_46 sp119_46 sp120_46 11.551961
Rsn119_46 sn119_46 sn120_46 11.551961
Rsp119_47 sp119_47 sp120_47 11.551961
Rsn119_47 sn119_47 sn120_47 11.551961
Rsp119_48 sp119_48 sp120_48 11.551961
Rsn119_48 sn119_48 sn120_48 11.551961
Rsp119_49 sp119_49 sp120_49 11.551961
Rsn119_49 sn119_49 sn120_49 11.551961
Rsp119_50 sp119_50 sp120_50 11.551961
Rsn119_50 sn119_50 sn120_50 11.551961
Rsp119_51 sp119_51 sp120_51 11.551961
Rsn119_51 sn119_51 sn120_51 11.551961
Rsp119_52 sp119_52 sp120_52 11.551961
Rsn119_52 sn119_52 sn120_52 11.551961
Rsp119_53 sp119_53 sp120_53 11.551961
Rsn119_53 sn119_53 sn120_53 11.551961
Rsp119_54 sp119_54 sp120_54 11.551961
Rsn119_54 sn119_54 sn120_54 11.551961
Rsp119_55 sp119_55 sp120_55 11.551961
Rsn119_55 sn119_55 sn120_55 11.551961
Rsp119_56 sp119_56 sp120_56 11.551961
Rsn119_56 sn119_56 sn120_56 11.551961
Rsp119_57 sp119_57 sp120_57 11.551961
Rsn119_57 sn119_57 sn120_57 11.551961
Rsp119_58 sp119_58 sp120_58 11.551961
Rsn119_58 sn119_58 sn120_58 11.551961
Rsp119_59 sp119_59 sp120_59 11.551961
Rsn119_59 sn119_59 sn120_59 11.551961
Rsp119_60 sp119_60 sp120_60 11.551961
Rsn119_60 sn119_60 sn120_60 11.551961
Rsp119_61 sp119_61 sp120_61 11.551961
Rsn119_61 sn119_61 sn120_61 11.551961
Rsp119_62 sp119_62 sp120_62 11.551961
Rsn119_62 sn119_62 sn120_62 11.551961
Rsp119_63 sp119_63 sp120_63 11.551961
Rsn119_63 sn119_63 sn120_63 11.551961
Rsp119_64 sp119_64 sp120_64 11.551961
Rsn119_64 sn119_64 sn120_64 11.551961
Rsp119_65 sp119_65 sp120_65 11.551961
Rsn119_65 sn119_65 sn120_65 11.551961
Rsp119_66 sp119_66 sp120_66 11.551961
Rsn119_66 sn119_66 sn120_66 11.551961
Rsp119_67 sp119_67 sp120_67 11.551961
Rsn119_67 sn119_67 sn120_67 11.551961
Rsp119_68 sp119_68 sp120_68 11.551961
Rsn119_68 sn119_68 sn120_68 11.551961
Rsp119_69 sp119_69 sp120_69 11.551961
Rsn119_69 sn119_69 sn120_69 11.551961
Rsp119_70 sp119_70 sp120_70 11.551961
Rsn119_70 sn119_70 sn120_70 11.551961
Rsp119_71 sp119_71 sp120_71 11.551961
Rsn119_71 sn119_71 sn120_71 11.551961
Rsp119_72 sp119_72 sp120_72 11.551961
Rsn119_72 sn119_72 sn120_72 11.551961
Rsp119_73 sp119_73 sp120_73 11.551961
Rsn119_73 sn119_73 sn120_73 11.551961
Rsp119_74 sp119_74 sp120_74 11.551961
Rsn119_74 sn119_74 sn120_74 11.551961
Rsp119_75 sp119_75 sp120_75 11.551961
Rsn119_75 sn119_75 sn120_75 11.551961
Rsp119_76 sp119_76 sp120_76 11.551961
Rsn119_76 sn119_76 sn120_76 11.551961
Rsp119_77 sp119_77 sp120_77 11.551961
Rsn119_77 sn119_77 sn120_77 11.551961
Rsp119_78 sp119_78 sp120_78 11.551961
Rsn119_78 sn119_78 sn120_78 11.551961
Rsp119_79 sp119_79 sp120_79 11.551961
Rsn119_79 sn119_79 sn120_79 11.551961
Rsp119_80 sp119_80 sp120_80 11.551961
Rsn119_80 sn119_80 sn120_80 11.551961
Rsp119_81 sp119_81 sp120_81 11.551961
Rsn119_81 sn119_81 sn120_81 11.551961
Rsp119_82 sp119_82 sp120_82 11.551961
Rsn119_82 sn119_82 sn120_82 11.551961
Rsp119_83 sp119_83 sp120_83 11.551961
Rsn119_83 sn119_83 sn120_83 11.551961
Rsp119_84 sp119_84 sp120_84 11.551961
Rsn119_84 sn119_84 sn120_84 11.551961
Rsp120_1 sp120_1 sp121_1 11.551961
Rsn120_1 sn120_1 sn121_1 11.551961
Rsp120_2 sp120_2 sp121_2 11.551961
Rsn120_2 sn120_2 sn121_2 11.551961
Rsp120_3 sp120_3 sp121_3 11.551961
Rsn120_3 sn120_3 sn121_3 11.551961
Rsp120_4 sp120_4 sp121_4 11.551961
Rsn120_4 sn120_4 sn121_4 11.551961
Rsp120_5 sp120_5 sp121_5 11.551961
Rsn120_5 sn120_5 sn121_5 11.551961
Rsp120_6 sp120_6 sp121_6 11.551961
Rsn120_6 sn120_6 sn121_6 11.551961
Rsp120_7 sp120_7 sp121_7 11.551961
Rsn120_7 sn120_7 sn121_7 11.551961
Rsp120_8 sp120_8 sp121_8 11.551961
Rsn120_8 sn120_8 sn121_8 11.551961
Rsp120_9 sp120_9 sp121_9 11.551961
Rsn120_9 sn120_9 sn121_9 11.551961
Rsp120_10 sp120_10 sp121_10 11.551961
Rsn120_10 sn120_10 sn121_10 11.551961
Rsp120_11 sp120_11 sp121_11 11.551961
Rsn120_11 sn120_11 sn121_11 11.551961
Rsp120_12 sp120_12 sp121_12 11.551961
Rsn120_12 sn120_12 sn121_12 11.551961
Rsp120_13 sp120_13 sp121_13 11.551961
Rsn120_13 sn120_13 sn121_13 11.551961
Rsp120_14 sp120_14 sp121_14 11.551961
Rsn120_14 sn120_14 sn121_14 11.551961
Rsp120_15 sp120_15 sp121_15 11.551961
Rsn120_15 sn120_15 sn121_15 11.551961
Rsp120_16 sp120_16 sp121_16 11.551961
Rsn120_16 sn120_16 sn121_16 11.551961
Rsp120_17 sp120_17 sp121_17 11.551961
Rsn120_17 sn120_17 sn121_17 11.551961
Rsp120_18 sp120_18 sp121_18 11.551961
Rsn120_18 sn120_18 sn121_18 11.551961
Rsp120_19 sp120_19 sp121_19 11.551961
Rsn120_19 sn120_19 sn121_19 11.551961
Rsp120_20 sp120_20 sp121_20 11.551961
Rsn120_20 sn120_20 sn121_20 11.551961
Rsp120_21 sp120_21 sp121_21 11.551961
Rsn120_21 sn120_21 sn121_21 11.551961
Rsp120_22 sp120_22 sp121_22 11.551961
Rsn120_22 sn120_22 sn121_22 11.551961
Rsp120_23 sp120_23 sp121_23 11.551961
Rsn120_23 sn120_23 sn121_23 11.551961
Rsp120_24 sp120_24 sp121_24 11.551961
Rsn120_24 sn120_24 sn121_24 11.551961
Rsp120_25 sp120_25 sp121_25 11.551961
Rsn120_25 sn120_25 sn121_25 11.551961
Rsp120_26 sp120_26 sp121_26 11.551961
Rsn120_26 sn120_26 sn121_26 11.551961
Rsp120_27 sp120_27 sp121_27 11.551961
Rsn120_27 sn120_27 sn121_27 11.551961
Rsp120_28 sp120_28 sp121_28 11.551961
Rsn120_28 sn120_28 sn121_28 11.551961
Rsp120_29 sp120_29 sp121_29 11.551961
Rsn120_29 sn120_29 sn121_29 11.551961
Rsp120_30 sp120_30 sp121_30 11.551961
Rsn120_30 sn120_30 sn121_30 11.551961
Rsp120_31 sp120_31 sp121_31 11.551961
Rsn120_31 sn120_31 sn121_31 11.551961
Rsp120_32 sp120_32 sp121_32 11.551961
Rsn120_32 sn120_32 sn121_32 11.551961
Rsp120_33 sp120_33 sp121_33 11.551961
Rsn120_33 sn120_33 sn121_33 11.551961
Rsp120_34 sp120_34 sp121_34 11.551961
Rsn120_34 sn120_34 sn121_34 11.551961
Rsp120_35 sp120_35 sp121_35 11.551961
Rsn120_35 sn120_35 sn121_35 11.551961
Rsp120_36 sp120_36 sp121_36 11.551961
Rsn120_36 sn120_36 sn121_36 11.551961
Rsp120_37 sp120_37 sp121_37 11.551961
Rsn120_37 sn120_37 sn121_37 11.551961
Rsp120_38 sp120_38 sp121_38 11.551961
Rsn120_38 sn120_38 sn121_38 11.551961
Rsp120_39 sp120_39 sp121_39 11.551961
Rsn120_39 sn120_39 sn121_39 11.551961
Rsp120_40 sp120_40 sp121_40 11.551961
Rsn120_40 sn120_40 sn121_40 11.551961
Rsp120_41 sp120_41 sp121_41 11.551961
Rsn120_41 sn120_41 sn121_41 11.551961
Rsp120_42 sp120_42 sp121_42 11.551961
Rsn120_42 sn120_42 sn121_42 11.551961
Rsp120_43 sp120_43 sp121_43 11.551961
Rsn120_43 sn120_43 sn121_43 11.551961
Rsp120_44 sp120_44 sp121_44 11.551961
Rsn120_44 sn120_44 sn121_44 11.551961
Rsp120_45 sp120_45 sp121_45 11.551961
Rsn120_45 sn120_45 sn121_45 11.551961
Rsp120_46 sp120_46 sp121_46 11.551961
Rsn120_46 sn120_46 sn121_46 11.551961
Rsp120_47 sp120_47 sp121_47 11.551961
Rsn120_47 sn120_47 sn121_47 11.551961
Rsp120_48 sp120_48 sp121_48 11.551961
Rsn120_48 sn120_48 sn121_48 11.551961
Rsp120_49 sp120_49 sp121_49 11.551961
Rsn120_49 sn120_49 sn121_49 11.551961
Rsp120_50 sp120_50 sp121_50 11.551961
Rsn120_50 sn120_50 sn121_50 11.551961
Rsp120_51 sp120_51 sp121_51 11.551961
Rsn120_51 sn120_51 sn121_51 11.551961
Rsp120_52 sp120_52 sp121_52 11.551961
Rsn120_52 sn120_52 sn121_52 11.551961
Rsp120_53 sp120_53 sp121_53 11.551961
Rsn120_53 sn120_53 sn121_53 11.551961
Rsp120_54 sp120_54 sp121_54 11.551961
Rsn120_54 sn120_54 sn121_54 11.551961
Rsp120_55 sp120_55 sp121_55 11.551961
Rsn120_55 sn120_55 sn121_55 11.551961
Rsp120_56 sp120_56 sp121_56 11.551961
Rsn120_56 sn120_56 sn121_56 11.551961
Rsp120_57 sp120_57 sp121_57 11.551961
Rsn120_57 sn120_57 sn121_57 11.551961
Rsp120_58 sp120_58 sp121_58 11.551961
Rsn120_58 sn120_58 sn121_58 11.551961
Rsp120_59 sp120_59 sp121_59 11.551961
Rsn120_59 sn120_59 sn121_59 11.551961
Rsp120_60 sp120_60 sp121_60 11.551961
Rsn120_60 sn120_60 sn121_60 11.551961
Rsp120_61 sp120_61 sp121_61 11.551961
Rsn120_61 sn120_61 sn121_61 11.551961
Rsp120_62 sp120_62 sp121_62 11.551961
Rsn120_62 sn120_62 sn121_62 11.551961
Rsp120_63 sp120_63 sp121_63 11.551961
Rsn120_63 sn120_63 sn121_63 11.551961
Rsp120_64 sp120_64 sp121_64 11.551961
Rsn120_64 sn120_64 sn121_64 11.551961
Rsp120_65 sp120_65 sp121_65 11.551961
Rsn120_65 sn120_65 sn121_65 11.551961
Rsp120_66 sp120_66 sp121_66 11.551961
Rsn120_66 sn120_66 sn121_66 11.551961
Rsp120_67 sp120_67 sp121_67 11.551961
Rsn120_67 sn120_67 sn121_67 11.551961
Rsp120_68 sp120_68 sp121_68 11.551961
Rsn120_68 sn120_68 sn121_68 11.551961
Rsp120_69 sp120_69 sp121_69 11.551961
Rsn120_69 sn120_69 sn121_69 11.551961
Rsp120_70 sp120_70 sp121_70 11.551961
Rsn120_70 sn120_70 sn121_70 11.551961
Rsp120_71 sp120_71 sp121_71 11.551961
Rsn120_71 sn120_71 sn121_71 11.551961
Rsp120_72 sp120_72 sp121_72 11.551961
Rsn120_72 sn120_72 sn121_72 11.551961
Rsp120_73 sp120_73 sp121_73 11.551961
Rsn120_73 sn120_73 sn121_73 11.551961
Rsp120_74 sp120_74 sp121_74 11.551961
Rsn120_74 sn120_74 sn121_74 11.551961
Rsp120_75 sp120_75 sp121_75 11.551961
Rsn120_75 sn120_75 sn121_75 11.551961
Rsp120_76 sp120_76 sp121_76 11.551961
Rsn120_76 sn120_76 sn121_76 11.551961
Rsp120_77 sp120_77 sp121_77 11.551961
Rsn120_77 sn120_77 sn121_77 11.551961
Rsp120_78 sp120_78 sp121_78 11.551961
Rsn120_78 sn120_78 sn121_78 11.551961
Rsp120_79 sp120_79 sp121_79 11.551961
Rsn120_79 sn120_79 sn121_79 11.551961
Rsp120_80 sp120_80 sp121_80 11.551961
Rsn120_80 sn120_80 sn121_80 11.551961
Rsp120_81 sp120_81 sp121_81 11.551961
Rsn120_81 sn120_81 sn121_81 11.551961
Rsp120_82 sp120_82 sp121_82 11.551961
Rsn120_82 sn120_82 sn121_82 11.551961
Rsp120_83 sp120_83 sp121_83 11.551961
Rsn120_83 sn120_83 sn121_83 11.551961
Rsp120_84 sp120_84 sp121_84 11.551961
Rsn120_84 sn120_84 sn121_84 11.551961
Rsp121_1 sp121_1 sp1_p4 11.551961
Rsn121_1 sn121_1 sn1_p4 11.551961
Rsp121_2 sp121_2 sp2_p4 11.551961
Rsn121_2 sn121_2 sn2_p4 11.551961
Rsp121_3 sp121_3 sp3_p4 11.551961
Rsn121_3 sn121_3 sn3_p4 11.551961
Rsp121_4 sp121_4 sp4_p4 11.551961
Rsn121_4 sn121_4 sn4_p4 11.551961
Rsp121_5 sp121_5 sp5_p4 11.551961
Rsn121_5 sn121_5 sn5_p4 11.551961
Rsp121_6 sp121_6 sp6_p4 11.551961
Rsn121_6 sn121_6 sn6_p4 11.551961
Rsp121_7 sp121_7 sp7_p4 11.551961
Rsn121_7 sn121_7 sn7_p4 11.551961
Rsp121_8 sp121_8 sp8_p4 11.551961
Rsn121_8 sn121_8 sn8_p4 11.551961
Rsp121_9 sp121_9 sp9_p4 11.551961
Rsn121_9 sn121_9 sn9_p4 11.551961
Rsp121_10 sp121_10 sp10_p4 11.551961
Rsn121_10 sn121_10 sn10_p4 11.551961
Rsp121_11 sp121_11 sp11_p4 11.551961
Rsn121_11 sn121_11 sn11_p4 11.551961
Rsp121_12 sp121_12 sp12_p4 11.551961
Rsn121_12 sn121_12 sn12_p4 11.551961
Rsp121_13 sp121_13 sp13_p4 11.551961
Rsn121_13 sn121_13 sn13_p4 11.551961
Rsp121_14 sp121_14 sp14_p4 11.551961
Rsn121_14 sn121_14 sn14_p4 11.551961
Rsp121_15 sp121_15 sp15_p4 11.551961
Rsn121_15 sn121_15 sn15_p4 11.551961
Rsp121_16 sp121_16 sp16_p4 11.551961
Rsn121_16 sn121_16 sn16_p4 11.551961
Rsp121_17 sp121_17 sp17_p4 11.551961
Rsn121_17 sn121_17 sn17_p4 11.551961
Rsp121_18 sp121_18 sp18_p4 11.551961
Rsn121_18 sn121_18 sn18_p4 11.551961
Rsp121_19 sp121_19 sp19_p4 11.551961
Rsn121_19 sn121_19 sn19_p4 11.551961
Rsp121_20 sp121_20 sp20_p4 11.551961
Rsn121_20 sn121_20 sn20_p4 11.551961
Rsp121_21 sp121_21 sp21_p4 11.551961
Rsn121_21 sn121_21 sn21_p4 11.551961
Rsp121_22 sp121_22 sp22_p4 11.551961
Rsn121_22 sn121_22 sn22_p4 11.551961
Rsp121_23 sp121_23 sp23_p4 11.551961
Rsn121_23 sn121_23 sn23_p4 11.551961
Rsp121_24 sp121_24 sp24_p4 11.551961
Rsn121_24 sn121_24 sn24_p4 11.551961
Rsp121_25 sp121_25 sp25_p4 11.551961
Rsn121_25 sn121_25 sn25_p4 11.551961
Rsp121_26 sp121_26 sp26_p4 11.551961
Rsn121_26 sn121_26 sn26_p4 11.551961
Rsp121_27 sp121_27 sp27_p4 11.551961
Rsn121_27 sn121_27 sn27_p4 11.551961
Rsp121_28 sp121_28 sp28_p4 11.551961
Rsn121_28 sn121_28 sn28_p4 11.551961
Rsp121_29 sp121_29 sp29_p4 11.551961
Rsn121_29 sn121_29 sn29_p4 11.551961
Rsp121_30 sp121_30 sp30_p4 11.551961
Rsn121_30 sn121_30 sn30_p4 11.551961
Rsp121_31 sp121_31 sp31_p4 11.551961
Rsn121_31 sn121_31 sn31_p4 11.551961
Rsp121_32 sp121_32 sp32_p4 11.551961
Rsn121_32 sn121_32 sn32_p4 11.551961
Rsp121_33 sp121_33 sp33_p4 11.551961
Rsn121_33 sn121_33 sn33_p4 11.551961
Rsp121_34 sp121_34 sp34_p4 11.551961
Rsn121_34 sn121_34 sn34_p4 11.551961
Rsp121_35 sp121_35 sp35_p4 11.551961
Rsn121_35 sn121_35 sn35_p4 11.551961
Rsp121_36 sp121_36 sp36_p4 11.551961
Rsn121_36 sn121_36 sn36_p4 11.551961
Rsp121_37 sp121_37 sp37_p4 11.551961
Rsn121_37 sn121_37 sn37_p4 11.551961
Rsp121_38 sp121_38 sp38_p4 11.551961
Rsn121_38 sn121_38 sn38_p4 11.551961
Rsp121_39 sp121_39 sp39_p4 11.551961
Rsn121_39 sn121_39 sn39_p4 11.551961
Rsp121_40 sp121_40 sp40_p4 11.551961
Rsn121_40 sn121_40 sn40_p4 11.551961
Rsp121_41 sp121_41 sp41_p4 11.551961
Rsn121_41 sn121_41 sn41_p4 11.551961
Rsp121_42 sp121_42 sp42_p4 11.551961
Rsn121_42 sn121_42 sn42_p4 11.551961
Rsp121_43 sp121_43 sp43_p4 11.551961
Rsn121_43 sn121_43 sn43_p4 11.551961
Rsp121_44 sp121_44 sp44_p4 11.551961
Rsn121_44 sn121_44 sn44_p4 11.551961
Rsp121_45 sp121_45 sp45_p4 11.551961
Rsn121_45 sn121_45 sn45_p4 11.551961
Rsp121_46 sp121_46 sp46_p4 11.551961
Rsn121_46 sn121_46 sn46_p4 11.551961
Rsp121_47 sp121_47 sp47_p4 11.551961
Rsn121_47 sn121_47 sn47_p4 11.551961
Rsp121_48 sp121_48 sp48_p4 11.551961
Rsn121_48 sn121_48 sn48_p4 11.551961
Rsp121_49 sp121_49 sp49_p4 11.551961
Rsn121_49 sn121_49 sn49_p4 11.551961
Rsp121_50 sp121_50 sp50_p4 11.551961
Rsn121_50 sn121_50 sn50_p4 11.551961
Rsp121_51 sp121_51 sp51_p4 11.551961
Rsn121_51 sn121_51 sn51_p4 11.551961
Rsp121_52 sp121_52 sp52_p4 11.551961
Rsn121_52 sn121_52 sn52_p4 11.551961
Rsp121_53 sp121_53 sp53_p4 11.551961
Rsn121_53 sn121_53 sn53_p4 11.551961
Rsp121_54 sp121_54 sp54_p4 11.551961
Rsn121_54 sn121_54 sn54_p4 11.551961
Rsp121_55 sp121_55 sp55_p4 11.551961
Rsn121_55 sn121_55 sn55_p4 11.551961
Rsp121_56 sp121_56 sp56_p4 11.551961
Rsn121_56 sn121_56 sn56_p4 11.551961
Rsp121_57 sp121_57 sp57_p4 11.551961
Rsn121_57 sn121_57 sn57_p4 11.551961
Rsp121_58 sp121_58 sp58_p4 11.551961
Rsn121_58 sn121_58 sn58_p4 11.551961
Rsp121_59 sp121_59 sp59_p4 11.551961
Rsn121_59 sn121_59 sn59_p4 11.551961
Rsp121_60 sp121_60 sp60_p4 11.551961
Rsn121_60 sn121_60 sn60_p4 11.551961
Rsp121_61 sp121_61 sp61_p4 11.551961
Rsn121_61 sn121_61 sn61_p4 11.551961
Rsp121_62 sp121_62 sp62_p4 11.551961
Rsn121_62 sn121_62 sn62_p4 11.551961
Rsp121_63 sp121_63 sp63_p4 11.551961
Rsn121_63 sn121_63 sn63_p4 11.551961
Rsp121_64 sp121_64 sp64_p4 11.551961
Rsn121_64 sn121_64 sn64_p4 11.551961
Rsp121_65 sp121_65 sp65_p4 11.551961
Rsn121_65 sn121_65 sn65_p4 11.551961
Rsp121_66 sp121_66 sp66_p4 11.551961
Rsn121_66 sn121_66 sn66_p4 11.551961
Rsp121_67 sp121_67 sp67_p4 11.551961
Rsn121_67 sn121_67 sn67_p4 11.551961
Rsp121_68 sp121_68 sp68_p4 11.551961
Rsn121_68 sn121_68 sn68_p4 11.551961
Rsp121_69 sp121_69 sp69_p4 11.551961
Rsn121_69 sn121_69 sn69_p4 11.551961
Rsp121_70 sp121_70 sp70_p4 11.551961
Rsn121_70 sn121_70 sn70_p4 11.551961
Rsp121_71 sp121_71 sp71_p4 11.551961
Rsn121_71 sn121_71 sn71_p4 11.551961
Rsp121_72 sp121_72 sp72_p4 11.551961
Rsn121_72 sn121_72 sn72_p4 11.551961
Rsp121_73 sp121_73 sp73_p4 11.551961
Rsn121_73 sn121_73 sn73_p4 11.551961
Rsp121_74 sp121_74 sp74_p4 11.551961
Rsn121_74 sn121_74 sn74_p4 11.551961
Rsp121_75 sp121_75 sp75_p4 11.551961
Rsn121_75 sn121_75 sn75_p4 11.551961
Rsp121_76 sp121_76 sp76_p4 11.551961
Rsn121_76 sn121_76 sn76_p4 11.551961
Rsp121_77 sp121_77 sp77_p4 11.551961
Rsn121_77 sn121_77 sn77_p4 11.551961
Rsp121_78 sp121_78 sp78_p4 11.551961
Rsn121_78 sn121_78 sn78_p4 11.551961
Rsp121_79 sp121_79 sp79_p4 11.551961
Rsn121_79 sn121_79 sn79_p4 11.551961
Rsp121_80 sp121_80 sp80_p4 11.551961
Rsn121_80 sn121_80 sn80_p4 11.551961
Rsp121_81 sp121_81 sp81_p4 11.551961
Rsn121_81 sn121_81 sn81_p4 11.551961
Rsp121_82 sp121_82 sp82_p4 11.551961
Rsn121_82 sn121_82 sn82_p4 11.551961
Rsp121_83 sp121_83 sp83_p4 11.551961
Rsn121_83 sn121_83 sn83_p4 11.551961
Rsp121_84 sp121_84 sp84_p4 11.551961
Rsn121_84 sn121_84 sn84_p4 11.551961


**********Weight Differntial Op-AMPS and Connecting Resistors****************

XDIFFw1_p1 sp1_p1 sn1_p1 nin1_1 diff2
Rconn1_p1 nin1_1 nin1 1m
XDIFFw2_p1 sp2_p1 sn2_p1 nin2_1 diff2
Rconn2_p1 nin2_1 nin2 1m
XDIFFw3_p1 sp3_p1 sn3_p1 nin3_1 diff2
Rconn3_p1 nin3_1 nin3 1m
XDIFFw4_p1 sp4_p1 sn4_p1 nin4_1 diff2
Rconn4_p1 nin4_1 nin4 1m
XDIFFw5_p1 sp5_p1 sn5_p1 nin5_1 diff2
Rconn5_p1 nin5_1 nin5 1m
XDIFFw6_p1 sp6_p1 sn6_p1 nin6_1 diff2
Rconn6_p1 nin6_1 nin6 1m
XDIFFw7_p1 sp7_p1 sn7_p1 nin7_1 diff2
Rconn7_p1 nin7_1 nin7 1m
XDIFFw8_p1 sp8_p1 sn8_p1 nin8_1 diff2
Rconn8_p1 nin8_1 nin8 1m
XDIFFw9_p1 sp9_p1 sn9_p1 nin9_1 diff2
Rconn9_p1 nin9_1 nin9 1m
XDIFFw10_p1 sp10_p1 sn10_p1 nin10_1 diff2
Rconn10_p1 nin10_1 nin10 1m
XDIFFw11_p1 sp11_p1 sn11_p1 nin11_1 diff2
Rconn11_p1 nin11_1 nin11 1m
XDIFFw12_p1 sp12_p1 sn12_p1 nin12_1 diff2
Rconn12_p1 nin12_1 nin12 1m
XDIFFw13_p1 sp13_p1 sn13_p1 nin13_1 diff2
Rconn13_p1 nin13_1 nin13 1m
XDIFFw14_p1 sp14_p1 sn14_p1 nin14_1 diff2
Rconn14_p1 nin14_1 nin14 1m
XDIFFw15_p1 sp15_p1 sn15_p1 nin15_1 diff2
Rconn15_p1 nin15_1 nin15 1m
XDIFFw16_p1 sp16_p1 sn16_p1 nin16_1 diff2
Rconn16_p1 nin16_1 nin16 1m
XDIFFw17_p1 sp17_p1 sn17_p1 nin17_1 diff2
Rconn17_p1 nin17_1 nin17 1m
XDIFFw18_p1 sp18_p1 sn18_p1 nin18_1 diff2
Rconn18_p1 nin18_1 nin18 1m
XDIFFw19_p1 sp19_p1 sn19_p1 nin19_1 diff2
Rconn19_p1 nin19_1 nin19 1m
XDIFFw20_p1 sp20_p1 sn20_p1 nin20_1 diff2
Rconn20_p1 nin20_1 nin20 1m
XDIFFw21_p1 sp21_p1 sn21_p1 nin21_1 diff2
Rconn21_p1 nin21_1 nin21 1m
XDIFFw22_p1 sp22_p1 sn22_p1 nin22_1 diff2
Rconn22_p1 nin22_1 nin22 1m
XDIFFw23_p1 sp23_p1 sn23_p1 nin23_1 diff2
Rconn23_p1 nin23_1 nin23 1m
XDIFFw24_p1 sp24_p1 sn24_p1 nin24_1 diff2
Rconn24_p1 nin24_1 nin24 1m
XDIFFw25_p1 sp25_p1 sn25_p1 nin25_1 diff2
Rconn25_p1 nin25_1 nin25 1m
XDIFFw26_p1 sp26_p1 sn26_p1 nin26_1 diff2
Rconn26_p1 nin26_1 nin26 1m
XDIFFw27_p1 sp27_p1 sn27_p1 nin27_1 diff2
Rconn27_p1 nin27_1 nin27 1m
XDIFFw28_p1 sp28_p1 sn28_p1 nin28_1 diff2
Rconn28_p1 nin28_1 nin28 1m
XDIFFw29_p1 sp29_p1 sn29_p1 nin29_1 diff2
Rconn29_p1 nin29_1 nin29 1m
XDIFFw30_p1 sp30_p1 sn30_p1 nin30_1 diff2
Rconn30_p1 nin30_1 nin30 1m
XDIFFw31_p1 sp31_p1 sn31_p1 nin31_1 diff2
Rconn31_p1 nin31_1 nin31 1m
XDIFFw32_p1 sp32_p1 sn32_p1 nin32_1 diff2
Rconn32_p1 nin32_1 nin32 1m
XDIFFw33_p1 sp33_p1 sn33_p1 nin33_1 diff2
Rconn33_p1 nin33_1 nin33 1m
XDIFFw34_p1 sp34_p1 sn34_p1 nin34_1 diff2
Rconn34_p1 nin34_1 nin34 1m
XDIFFw35_p1 sp35_p1 sn35_p1 nin35_1 diff2
Rconn35_p1 nin35_1 nin35 1m
XDIFFw36_p1 sp36_p1 sn36_p1 nin36_1 diff2
Rconn36_p1 nin36_1 nin36 1m
XDIFFw37_p1 sp37_p1 sn37_p1 nin37_1 diff2
Rconn37_p1 nin37_1 nin37 1m
XDIFFw38_p1 sp38_p1 sn38_p1 nin38_1 diff2
Rconn38_p1 nin38_1 nin38 1m
XDIFFw39_p1 sp39_p1 sn39_p1 nin39_1 diff2
Rconn39_p1 nin39_1 nin39 1m
XDIFFw40_p1 sp40_p1 sn40_p1 nin40_1 diff2
Rconn40_p1 nin40_1 nin40 1m
XDIFFw41_p1 sp41_p1 sn41_p1 nin41_1 diff2
Rconn41_p1 nin41_1 nin41 1m
XDIFFw42_p1 sp42_p1 sn42_p1 nin42_1 diff2
Rconn42_p1 nin42_1 nin42 1m
XDIFFw43_p1 sp43_p1 sn43_p1 nin43_1 diff2
Rconn43_p1 nin43_1 nin43 1m
XDIFFw44_p1 sp44_p1 sn44_p1 nin44_1 diff2
Rconn44_p1 nin44_1 nin44 1m
XDIFFw45_p1 sp45_p1 sn45_p1 nin45_1 diff2
Rconn45_p1 nin45_1 nin45 1m
XDIFFw46_p1 sp46_p1 sn46_p1 nin46_1 diff2
Rconn46_p1 nin46_1 nin46 1m
XDIFFw47_p1 sp47_p1 sn47_p1 nin47_1 diff2
Rconn47_p1 nin47_1 nin47 1m
XDIFFw48_p1 sp48_p1 sn48_p1 nin48_1 diff2
Rconn48_p1 nin48_1 nin48 1m
XDIFFw49_p1 sp49_p1 sn49_p1 nin49_1 diff2
Rconn49_p1 nin49_1 nin49 1m
XDIFFw50_p1 sp50_p1 sn50_p1 nin50_1 diff2
Rconn50_p1 nin50_1 nin50 1m
XDIFFw51_p1 sp51_p1 sn51_p1 nin51_1 diff2
Rconn51_p1 nin51_1 nin51 1m
XDIFFw52_p1 sp52_p1 sn52_p1 nin52_1 diff2
Rconn52_p1 nin52_1 nin52 1m
XDIFFw53_p1 sp53_p1 sn53_p1 nin53_1 diff2
Rconn53_p1 nin53_1 nin53 1m
XDIFFw54_p1 sp54_p1 sn54_p1 nin54_1 diff2
Rconn54_p1 nin54_1 nin54 1m
XDIFFw55_p1 sp55_p1 sn55_p1 nin55_1 diff2
Rconn55_p1 nin55_1 nin55 1m
XDIFFw56_p1 sp56_p1 sn56_p1 nin56_1 diff2
Rconn56_p1 nin56_1 nin56 1m
XDIFFw57_p1 sp57_p1 sn57_p1 nin57_1 diff2
Rconn57_p1 nin57_1 nin57 1m
XDIFFw58_p1 sp58_p1 sn58_p1 nin58_1 diff2
Rconn58_p1 nin58_1 nin58 1m
XDIFFw59_p1 sp59_p1 sn59_p1 nin59_1 diff2
Rconn59_p1 nin59_1 nin59 1m
XDIFFw60_p1 sp60_p1 sn60_p1 nin60_1 diff2
Rconn60_p1 nin60_1 nin60 1m
XDIFFw61_p1 sp61_p1 sn61_p1 nin61_1 diff2
Rconn61_p1 nin61_1 nin61 1m
XDIFFw62_p1 sp62_p1 sn62_p1 nin62_1 diff2
Rconn62_p1 nin62_1 nin62 1m
XDIFFw63_p1 sp63_p1 sn63_p1 nin63_1 diff2
Rconn63_p1 nin63_1 nin63 1m
XDIFFw64_p1 sp64_p1 sn64_p1 nin64_1 diff2
Rconn64_p1 nin64_1 nin64 1m
XDIFFw65_p1 sp65_p1 sn65_p1 nin65_1 diff2
Rconn65_p1 nin65_1 nin65 1m
XDIFFw66_p1 sp66_p1 sn66_p1 nin66_1 diff2
Rconn66_p1 nin66_1 nin66 1m
XDIFFw67_p1 sp67_p1 sn67_p1 nin67_1 diff2
Rconn67_p1 nin67_1 nin67 1m
XDIFFw68_p1 sp68_p1 sn68_p1 nin68_1 diff2
Rconn68_p1 nin68_1 nin68 1m
XDIFFw69_p1 sp69_p1 sn69_p1 nin69_1 diff2
Rconn69_p1 nin69_1 nin69 1m
XDIFFw70_p1 sp70_p1 sn70_p1 nin70_1 diff2
Rconn70_p1 nin70_1 nin70 1m
XDIFFw71_p1 sp71_p1 sn71_p1 nin71_1 diff2
Rconn71_p1 nin71_1 nin71 1m
XDIFFw72_p1 sp72_p1 sn72_p1 nin72_1 diff2
Rconn72_p1 nin72_1 nin72 1m
XDIFFw73_p1 sp73_p1 sn73_p1 nin73_1 diff2
Rconn73_p1 nin73_1 nin73 1m
XDIFFw74_p1 sp74_p1 sn74_p1 nin74_1 diff2
Rconn74_p1 nin74_1 nin74 1m
XDIFFw75_p1 sp75_p1 sn75_p1 nin75_1 diff2
Rconn75_p1 nin75_1 nin75 1m
XDIFFw76_p1 sp76_p1 sn76_p1 nin76_1 diff2
Rconn76_p1 nin76_1 nin76 1m
XDIFFw77_p1 sp77_p1 sn77_p1 nin77_1 diff2
Rconn77_p1 nin77_1 nin77 1m
XDIFFw78_p1 sp78_p1 sn78_p1 nin78_1 diff2
Rconn78_p1 nin78_1 nin78 1m
XDIFFw79_p1 sp79_p1 sn79_p1 nin79_1 diff2
Rconn79_p1 nin79_1 nin79 1m
XDIFFw80_p1 sp80_p1 sn80_p1 nin80_1 diff2
Rconn80_p1 nin80_1 nin80 1m
XDIFFw81_p1 sp81_p1 sn81_p1 nin81_1 diff2
Rconn81_p1 nin81_1 nin81 1m
XDIFFw82_p1 sp82_p1 sn82_p1 nin82_1 diff2
Rconn82_p1 nin82_1 nin82 1m
XDIFFw83_p1 sp83_p1 sn83_p1 nin83_1 diff2
Rconn83_p1 nin83_1 nin83 1m
XDIFFw84_p1 sp84_p1 sn84_p1 nin84_1 diff2
Rconn84_p1 nin84_1 nin84 1m
XDIFFw1_p2 sp1_p2 sn1_p2 nin1_2 diff2
Rconn1_p2 nin1_2 nin1 1m
XDIFFw2_p2 sp2_p2 sn2_p2 nin2_2 diff2
Rconn2_p2 nin2_2 nin2 1m
XDIFFw3_p2 sp3_p2 sn3_p2 nin3_2 diff2
Rconn3_p2 nin3_2 nin3 1m
XDIFFw4_p2 sp4_p2 sn4_p2 nin4_2 diff2
Rconn4_p2 nin4_2 nin4 1m
XDIFFw5_p2 sp5_p2 sn5_p2 nin5_2 diff2
Rconn5_p2 nin5_2 nin5 1m
XDIFFw6_p2 sp6_p2 sn6_p2 nin6_2 diff2
Rconn6_p2 nin6_2 nin6 1m
XDIFFw7_p2 sp7_p2 sn7_p2 nin7_2 diff2
Rconn7_p2 nin7_2 nin7 1m
XDIFFw8_p2 sp8_p2 sn8_p2 nin8_2 diff2
Rconn8_p2 nin8_2 nin8 1m
XDIFFw9_p2 sp9_p2 sn9_p2 nin9_2 diff2
Rconn9_p2 nin9_2 nin9 1m
XDIFFw10_p2 sp10_p2 sn10_p2 nin10_2 diff2
Rconn10_p2 nin10_2 nin10 1m
XDIFFw11_p2 sp11_p2 sn11_p2 nin11_2 diff2
Rconn11_p2 nin11_2 nin11 1m
XDIFFw12_p2 sp12_p2 sn12_p2 nin12_2 diff2
Rconn12_p2 nin12_2 nin12 1m
XDIFFw13_p2 sp13_p2 sn13_p2 nin13_2 diff2
Rconn13_p2 nin13_2 nin13 1m
XDIFFw14_p2 sp14_p2 sn14_p2 nin14_2 diff2
Rconn14_p2 nin14_2 nin14 1m
XDIFFw15_p2 sp15_p2 sn15_p2 nin15_2 diff2
Rconn15_p2 nin15_2 nin15 1m
XDIFFw16_p2 sp16_p2 sn16_p2 nin16_2 diff2
Rconn16_p2 nin16_2 nin16 1m
XDIFFw17_p2 sp17_p2 sn17_p2 nin17_2 diff2
Rconn17_p2 nin17_2 nin17 1m
XDIFFw18_p2 sp18_p2 sn18_p2 nin18_2 diff2
Rconn18_p2 nin18_2 nin18 1m
XDIFFw19_p2 sp19_p2 sn19_p2 nin19_2 diff2
Rconn19_p2 nin19_2 nin19 1m
XDIFFw20_p2 sp20_p2 sn20_p2 nin20_2 diff2
Rconn20_p2 nin20_2 nin20 1m
XDIFFw21_p2 sp21_p2 sn21_p2 nin21_2 diff2
Rconn21_p2 nin21_2 nin21 1m
XDIFFw22_p2 sp22_p2 sn22_p2 nin22_2 diff2
Rconn22_p2 nin22_2 nin22 1m
XDIFFw23_p2 sp23_p2 sn23_p2 nin23_2 diff2
Rconn23_p2 nin23_2 nin23 1m
XDIFFw24_p2 sp24_p2 sn24_p2 nin24_2 diff2
Rconn24_p2 nin24_2 nin24 1m
XDIFFw25_p2 sp25_p2 sn25_p2 nin25_2 diff2
Rconn25_p2 nin25_2 nin25 1m
XDIFFw26_p2 sp26_p2 sn26_p2 nin26_2 diff2
Rconn26_p2 nin26_2 nin26 1m
XDIFFw27_p2 sp27_p2 sn27_p2 nin27_2 diff2
Rconn27_p2 nin27_2 nin27 1m
XDIFFw28_p2 sp28_p2 sn28_p2 nin28_2 diff2
Rconn28_p2 nin28_2 nin28 1m
XDIFFw29_p2 sp29_p2 sn29_p2 nin29_2 diff2
Rconn29_p2 nin29_2 nin29 1m
XDIFFw30_p2 sp30_p2 sn30_p2 nin30_2 diff2
Rconn30_p2 nin30_2 nin30 1m
XDIFFw31_p2 sp31_p2 sn31_p2 nin31_2 diff2
Rconn31_p2 nin31_2 nin31 1m
XDIFFw32_p2 sp32_p2 sn32_p2 nin32_2 diff2
Rconn32_p2 nin32_2 nin32 1m
XDIFFw33_p2 sp33_p2 sn33_p2 nin33_2 diff2
Rconn33_p2 nin33_2 nin33 1m
XDIFFw34_p2 sp34_p2 sn34_p2 nin34_2 diff2
Rconn34_p2 nin34_2 nin34 1m
XDIFFw35_p2 sp35_p2 sn35_p2 nin35_2 diff2
Rconn35_p2 nin35_2 nin35 1m
XDIFFw36_p2 sp36_p2 sn36_p2 nin36_2 diff2
Rconn36_p2 nin36_2 nin36 1m
XDIFFw37_p2 sp37_p2 sn37_p2 nin37_2 diff2
Rconn37_p2 nin37_2 nin37 1m
XDIFFw38_p2 sp38_p2 sn38_p2 nin38_2 diff2
Rconn38_p2 nin38_2 nin38 1m
XDIFFw39_p2 sp39_p2 sn39_p2 nin39_2 diff2
Rconn39_p2 nin39_2 nin39 1m
XDIFFw40_p2 sp40_p2 sn40_p2 nin40_2 diff2
Rconn40_p2 nin40_2 nin40 1m
XDIFFw41_p2 sp41_p2 sn41_p2 nin41_2 diff2
Rconn41_p2 nin41_2 nin41 1m
XDIFFw42_p2 sp42_p2 sn42_p2 nin42_2 diff2
Rconn42_p2 nin42_2 nin42 1m
XDIFFw43_p2 sp43_p2 sn43_p2 nin43_2 diff2
Rconn43_p2 nin43_2 nin43 1m
XDIFFw44_p2 sp44_p2 sn44_p2 nin44_2 diff2
Rconn44_p2 nin44_2 nin44 1m
XDIFFw45_p2 sp45_p2 sn45_p2 nin45_2 diff2
Rconn45_p2 nin45_2 nin45 1m
XDIFFw46_p2 sp46_p2 sn46_p2 nin46_2 diff2
Rconn46_p2 nin46_2 nin46 1m
XDIFFw47_p2 sp47_p2 sn47_p2 nin47_2 diff2
Rconn47_p2 nin47_2 nin47 1m
XDIFFw48_p2 sp48_p2 sn48_p2 nin48_2 diff2
Rconn48_p2 nin48_2 nin48 1m
XDIFFw49_p2 sp49_p2 sn49_p2 nin49_2 diff2
Rconn49_p2 nin49_2 nin49 1m
XDIFFw50_p2 sp50_p2 sn50_p2 nin50_2 diff2
Rconn50_p2 nin50_2 nin50 1m
XDIFFw51_p2 sp51_p2 sn51_p2 nin51_2 diff2
Rconn51_p2 nin51_2 nin51 1m
XDIFFw52_p2 sp52_p2 sn52_p2 nin52_2 diff2
Rconn52_p2 nin52_2 nin52 1m
XDIFFw53_p2 sp53_p2 sn53_p2 nin53_2 diff2
Rconn53_p2 nin53_2 nin53 1m
XDIFFw54_p2 sp54_p2 sn54_p2 nin54_2 diff2
Rconn54_p2 nin54_2 nin54 1m
XDIFFw55_p2 sp55_p2 sn55_p2 nin55_2 diff2
Rconn55_p2 nin55_2 nin55 1m
XDIFFw56_p2 sp56_p2 sn56_p2 nin56_2 diff2
Rconn56_p2 nin56_2 nin56 1m
XDIFFw57_p2 sp57_p2 sn57_p2 nin57_2 diff2
Rconn57_p2 nin57_2 nin57 1m
XDIFFw58_p2 sp58_p2 sn58_p2 nin58_2 diff2
Rconn58_p2 nin58_2 nin58 1m
XDIFFw59_p2 sp59_p2 sn59_p2 nin59_2 diff2
Rconn59_p2 nin59_2 nin59 1m
XDIFFw60_p2 sp60_p2 sn60_p2 nin60_2 diff2
Rconn60_p2 nin60_2 nin60 1m
XDIFFw61_p2 sp61_p2 sn61_p2 nin61_2 diff2
Rconn61_p2 nin61_2 nin61 1m
XDIFFw62_p2 sp62_p2 sn62_p2 nin62_2 diff2
Rconn62_p2 nin62_2 nin62 1m
XDIFFw63_p2 sp63_p2 sn63_p2 nin63_2 diff2
Rconn63_p2 nin63_2 nin63 1m
XDIFFw64_p2 sp64_p2 sn64_p2 nin64_2 diff2
Rconn64_p2 nin64_2 nin64 1m
XDIFFw65_p2 sp65_p2 sn65_p2 nin65_2 diff2
Rconn65_p2 nin65_2 nin65 1m
XDIFFw66_p2 sp66_p2 sn66_p2 nin66_2 diff2
Rconn66_p2 nin66_2 nin66 1m
XDIFFw67_p2 sp67_p2 sn67_p2 nin67_2 diff2
Rconn67_p2 nin67_2 nin67 1m
XDIFFw68_p2 sp68_p2 sn68_p2 nin68_2 diff2
Rconn68_p2 nin68_2 nin68 1m
XDIFFw69_p2 sp69_p2 sn69_p2 nin69_2 diff2
Rconn69_p2 nin69_2 nin69 1m
XDIFFw70_p2 sp70_p2 sn70_p2 nin70_2 diff2
Rconn70_p2 nin70_2 nin70 1m
XDIFFw71_p2 sp71_p2 sn71_p2 nin71_2 diff2
Rconn71_p2 nin71_2 nin71 1m
XDIFFw72_p2 sp72_p2 sn72_p2 nin72_2 diff2
Rconn72_p2 nin72_2 nin72 1m
XDIFFw73_p2 sp73_p2 sn73_p2 nin73_2 diff2
Rconn73_p2 nin73_2 nin73 1m
XDIFFw74_p2 sp74_p2 sn74_p2 nin74_2 diff2
Rconn74_p2 nin74_2 nin74 1m
XDIFFw75_p2 sp75_p2 sn75_p2 nin75_2 diff2
Rconn75_p2 nin75_2 nin75 1m
XDIFFw76_p2 sp76_p2 sn76_p2 nin76_2 diff2
Rconn76_p2 nin76_2 nin76 1m
XDIFFw77_p2 sp77_p2 sn77_p2 nin77_2 diff2
Rconn77_p2 nin77_2 nin77 1m
XDIFFw78_p2 sp78_p2 sn78_p2 nin78_2 diff2
Rconn78_p2 nin78_2 nin78 1m
XDIFFw79_p2 sp79_p2 sn79_p2 nin79_2 diff2
Rconn79_p2 nin79_2 nin79 1m
XDIFFw80_p2 sp80_p2 sn80_p2 nin80_2 diff2
Rconn80_p2 nin80_2 nin80 1m
XDIFFw81_p2 sp81_p2 sn81_p2 nin81_2 diff2
Rconn81_p2 nin81_2 nin81 1m
XDIFFw82_p2 sp82_p2 sn82_p2 nin82_2 diff2
Rconn82_p2 nin82_2 nin82 1m
XDIFFw83_p2 sp83_p2 sn83_p2 nin83_2 diff2
Rconn83_p2 nin83_2 nin83 1m
XDIFFw84_p2 sp84_p2 sn84_p2 nin84_2 diff2
Rconn84_p2 nin84_2 nin84 1m
XDIFFw1_p3 sp1_p3 sn1_p3 nin1_3 diff2
Rconn1_p3 nin1_3 nin1 1m
XDIFFw2_p3 sp2_p3 sn2_p3 nin2_3 diff2
Rconn2_p3 nin2_3 nin2 1m
XDIFFw3_p3 sp3_p3 sn3_p3 nin3_3 diff2
Rconn3_p3 nin3_3 nin3 1m
XDIFFw4_p3 sp4_p3 sn4_p3 nin4_3 diff2
Rconn4_p3 nin4_3 nin4 1m
XDIFFw5_p3 sp5_p3 sn5_p3 nin5_3 diff2
Rconn5_p3 nin5_3 nin5 1m
XDIFFw6_p3 sp6_p3 sn6_p3 nin6_3 diff2
Rconn6_p3 nin6_3 nin6 1m
XDIFFw7_p3 sp7_p3 sn7_p3 nin7_3 diff2
Rconn7_p3 nin7_3 nin7 1m
XDIFFw8_p3 sp8_p3 sn8_p3 nin8_3 diff2
Rconn8_p3 nin8_3 nin8 1m
XDIFFw9_p3 sp9_p3 sn9_p3 nin9_3 diff2
Rconn9_p3 nin9_3 nin9 1m
XDIFFw10_p3 sp10_p3 sn10_p3 nin10_3 diff2
Rconn10_p3 nin10_3 nin10 1m
XDIFFw11_p3 sp11_p3 sn11_p3 nin11_3 diff2
Rconn11_p3 nin11_3 nin11 1m
XDIFFw12_p3 sp12_p3 sn12_p3 nin12_3 diff2
Rconn12_p3 nin12_3 nin12 1m
XDIFFw13_p3 sp13_p3 sn13_p3 nin13_3 diff2
Rconn13_p3 nin13_3 nin13 1m
XDIFFw14_p3 sp14_p3 sn14_p3 nin14_3 diff2
Rconn14_p3 nin14_3 nin14 1m
XDIFFw15_p3 sp15_p3 sn15_p3 nin15_3 diff2
Rconn15_p3 nin15_3 nin15 1m
XDIFFw16_p3 sp16_p3 sn16_p3 nin16_3 diff2
Rconn16_p3 nin16_3 nin16 1m
XDIFFw17_p3 sp17_p3 sn17_p3 nin17_3 diff2
Rconn17_p3 nin17_3 nin17 1m
XDIFFw18_p3 sp18_p3 sn18_p3 nin18_3 diff2
Rconn18_p3 nin18_3 nin18 1m
XDIFFw19_p3 sp19_p3 sn19_p3 nin19_3 diff2
Rconn19_p3 nin19_3 nin19 1m
XDIFFw20_p3 sp20_p3 sn20_p3 nin20_3 diff2
Rconn20_p3 nin20_3 nin20 1m
XDIFFw21_p3 sp21_p3 sn21_p3 nin21_3 diff2
Rconn21_p3 nin21_3 nin21 1m
XDIFFw22_p3 sp22_p3 sn22_p3 nin22_3 diff2
Rconn22_p3 nin22_3 nin22 1m
XDIFFw23_p3 sp23_p3 sn23_p3 nin23_3 diff2
Rconn23_p3 nin23_3 nin23 1m
XDIFFw24_p3 sp24_p3 sn24_p3 nin24_3 diff2
Rconn24_p3 nin24_3 nin24 1m
XDIFFw25_p3 sp25_p3 sn25_p3 nin25_3 diff2
Rconn25_p3 nin25_3 nin25 1m
XDIFFw26_p3 sp26_p3 sn26_p3 nin26_3 diff2
Rconn26_p3 nin26_3 nin26 1m
XDIFFw27_p3 sp27_p3 sn27_p3 nin27_3 diff2
Rconn27_p3 nin27_3 nin27 1m
XDIFFw28_p3 sp28_p3 sn28_p3 nin28_3 diff2
Rconn28_p3 nin28_3 nin28 1m
XDIFFw29_p3 sp29_p3 sn29_p3 nin29_3 diff2
Rconn29_p3 nin29_3 nin29 1m
XDIFFw30_p3 sp30_p3 sn30_p3 nin30_3 diff2
Rconn30_p3 nin30_3 nin30 1m
XDIFFw31_p3 sp31_p3 sn31_p3 nin31_3 diff2
Rconn31_p3 nin31_3 nin31 1m
XDIFFw32_p3 sp32_p3 sn32_p3 nin32_3 diff2
Rconn32_p3 nin32_3 nin32 1m
XDIFFw33_p3 sp33_p3 sn33_p3 nin33_3 diff2
Rconn33_p3 nin33_3 nin33 1m
XDIFFw34_p3 sp34_p3 sn34_p3 nin34_3 diff2
Rconn34_p3 nin34_3 nin34 1m
XDIFFw35_p3 sp35_p3 sn35_p3 nin35_3 diff2
Rconn35_p3 nin35_3 nin35 1m
XDIFFw36_p3 sp36_p3 sn36_p3 nin36_3 diff2
Rconn36_p3 nin36_3 nin36 1m
XDIFFw37_p3 sp37_p3 sn37_p3 nin37_3 diff2
Rconn37_p3 nin37_3 nin37 1m
XDIFFw38_p3 sp38_p3 sn38_p3 nin38_3 diff2
Rconn38_p3 nin38_3 nin38 1m
XDIFFw39_p3 sp39_p3 sn39_p3 nin39_3 diff2
Rconn39_p3 nin39_3 nin39 1m
XDIFFw40_p3 sp40_p3 sn40_p3 nin40_3 diff2
Rconn40_p3 nin40_3 nin40 1m
XDIFFw41_p3 sp41_p3 sn41_p3 nin41_3 diff2
Rconn41_p3 nin41_3 nin41 1m
XDIFFw42_p3 sp42_p3 sn42_p3 nin42_3 diff2
Rconn42_p3 nin42_3 nin42 1m
XDIFFw43_p3 sp43_p3 sn43_p3 nin43_3 diff2
Rconn43_p3 nin43_3 nin43 1m
XDIFFw44_p3 sp44_p3 sn44_p3 nin44_3 diff2
Rconn44_p3 nin44_3 nin44 1m
XDIFFw45_p3 sp45_p3 sn45_p3 nin45_3 diff2
Rconn45_p3 nin45_3 nin45 1m
XDIFFw46_p3 sp46_p3 sn46_p3 nin46_3 diff2
Rconn46_p3 nin46_3 nin46 1m
XDIFFw47_p3 sp47_p3 sn47_p3 nin47_3 diff2
Rconn47_p3 nin47_3 nin47 1m
XDIFFw48_p3 sp48_p3 sn48_p3 nin48_3 diff2
Rconn48_p3 nin48_3 nin48 1m
XDIFFw49_p3 sp49_p3 sn49_p3 nin49_3 diff2
Rconn49_p3 nin49_3 nin49 1m
XDIFFw50_p3 sp50_p3 sn50_p3 nin50_3 diff2
Rconn50_p3 nin50_3 nin50 1m
XDIFFw51_p3 sp51_p3 sn51_p3 nin51_3 diff2
Rconn51_p3 nin51_3 nin51 1m
XDIFFw52_p3 sp52_p3 sn52_p3 nin52_3 diff2
Rconn52_p3 nin52_3 nin52 1m
XDIFFw53_p3 sp53_p3 sn53_p3 nin53_3 diff2
Rconn53_p3 nin53_3 nin53 1m
XDIFFw54_p3 sp54_p3 sn54_p3 nin54_3 diff2
Rconn54_p3 nin54_3 nin54 1m
XDIFFw55_p3 sp55_p3 sn55_p3 nin55_3 diff2
Rconn55_p3 nin55_3 nin55 1m
XDIFFw56_p3 sp56_p3 sn56_p3 nin56_3 diff2
Rconn56_p3 nin56_3 nin56 1m
XDIFFw57_p3 sp57_p3 sn57_p3 nin57_3 diff2
Rconn57_p3 nin57_3 nin57 1m
XDIFFw58_p3 sp58_p3 sn58_p3 nin58_3 diff2
Rconn58_p3 nin58_3 nin58 1m
XDIFFw59_p3 sp59_p3 sn59_p3 nin59_3 diff2
Rconn59_p3 nin59_3 nin59 1m
XDIFFw60_p3 sp60_p3 sn60_p3 nin60_3 diff2
Rconn60_p3 nin60_3 nin60 1m
XDIFFw61_p3 sp61_p3 sn61_p3 nin61_3 diff2
Rconn61_p3 nin61_3 nin61 1m
XDIFFw62_p3 sp62_p3 sn62_p3 nin62_3 diff2
Rconn62_p3 nin62_3 nin62 1m
XDIFFw63_p3 sp63_p3 sn63_p3 nin63_3 diff2
Rconn63_p3 nin63_3 nin63 1m
XDIFFw64_p3 sp64_p3 sn64_p3 nin64_3 diff2
Rconn64_p3 nin64_3 nin64 1m
XDIFFw65_p3 sp65_p3 sn65_p3 nin65_3 diff2
Rconn65_p3 nin65_3 nin65 1m
XDIFFw66_p3 sp66_p3 sn66_p3 nin66_3 diff2
Rconn66_p3 nin66_3 nin66 1m
XDIFFw67_p3 sp67_p3 sn67_p3 nin67_3 diff2
Rconn67_p3 nin67_3 nin67 1m
XDIFFw68_p3 sp68_p3 sn68_p3 nin68_3 diff2
Rconn68_p3 nin68_3 nin68 1m
XDIFFw69_p3 sp69_p3 sn69_p3 nin69_3 diff2
Rconn69_p3 nin69_3 nin69 1m
XDIFFw70_p3 sp70_p3 sn70_p3 nin70_3 diff2
Rconn70_p3 nin70_3 nin70 1m
XDIFFw71_p3 sp71_p3 sn71_p3 nin71_3 diff2
Rconn71_p3 nin71_3 nin71 1m
XDIFFw72_p3 sp72_p3 sn72_p3 nin72_3 diff2
Rconn72_p3 nin72_3 nin72 1m
XDIFFw73_p3 sp73_p3 sn73_p3 nin73_3 diff2
Rconn73_p3 nin73_3 nin73 1m
XDIFFw74_p3 sp74_p3 sn74_p3 nin74_3 diff2
Rconn74_p3 nin74_3 nin74 1m
XDIFFw75_p3 sp75_p3 sn75_p3 nin75_3 diff2
Rconn75_p3 nin75_3 nin75 1m
XDIFFw76_p3 sp76_p3 sn76_p3 nin76_3 diff2
Rconn76_p3 nin76_3 nin76 1m
XDIFFw77_p3 sp77_p3 sn77_p3 nin77_3 diff2
Rconn77_p3 nin77_3 nin77 1m
XDIFFw78_p3 sp78_p3 sn78_p3 nin78_3 diff2
Rconn78_p3 nin78_3 nin78 1m
XDIFFw79_p3 sp79_p3 sn79_p3 nin79_3 diff2
Rconn79_p3 nin79_3 nin79 1m
XDIFFw80_p3 sp80_p3 sn80_p3 nin80_3 diff2
Rconn80_p3 nin80_3 nin80 1m
XDIFFw81_p3 sp81_p3 sn81_p3 nin81_3 diff2
Rconn81_p3 nin81_3 nin81 1m
XDIFFw82_p3 sp82_p3 sn82_p3 nin82_3 diff2
Rconn82_p3 nin82_3 nin82 1m
XDIFFw83_p3 sp83_p3 sn83_p3 nin83_3 diff2
Rconn83_p3 nin83_3 nin83 1m
XDIFFw84_p3 sp84_p3 sn84_p3 nin84_3 diff2
Rconn84_p3 nin84_3 nin84 1m
XDIFFw1_p4 sp1_p4 sn1_p4 nin1_4 diff2
Rconn1_p4 nin1_4 nin1 1m
XDIFFw2_p4 sp2_p4 sn2_p4 nin2_4 diff2
Rconn2_p4 nin2_4 nin2 1m
XDIFFw3_p4 sp3_p4 sn3_p4 nin3_4 diff2
Rconn3_p4 nin3_4 nin3 1m
XDIFFw4_p4 sp4_p4 sn4_p4 nin4_4 diff2
Rconn4_p4 nin4_4 nin4 1m
XDIFFw5_p4 sp5_p4 sn5_p4 nin5_4 diff2
Rconn5_p4 nin5_4 nin5 1m
XDIFFw6_p4 sp6_p4 sn6_p4 nin6_4 diff2
Rconn6_p4 nin6_4 nin6 1m
XDIFFw7_p4 sp7_p4 sn7_p4 nin7_4 diff2
Rconn7_p4 nin7_4 nin7 1m
XDIFFw8_p4 sp8_p4 sn8_p4 nin8_4 diff2
Rconn8_p4 nin8_4 nin8 1m
XDIFFw9_p4 sp9_p4 sn9_p4 nin9_4 diff2
Rconn9_p4 nin9_4 nin9 1m
XDIFFw10_p4 sp10_p4 sn10_p4 nin10_4 diff2
Rconn10_p4 nin10_4 nin10 1m
XDIFFw11_p4 sp11_p4 sn11_p4 nin11_4 diff2
Rconn11_p4 nin11_4 nin11 1m
XDIFFw12_p4 sp12_p4 sn12_p4 nin12_4 diff2
Rconn12_p4 nin12_4 nin12 1m
XDIFFw13_p4 sp13_p4 sn13_p4 nin13_4 diff2
Rconn13_p4 nin13_4 nin13 1m
XDIFFw14_p4 sp14_p4 sn14_p4 nin14_4 diff2
Rconn14_p4 nin14_4 nin14 1m
XDIFFw15_p4 sp15_p4 sn15_p4 nin15_4 diff2
Rconn15_p4 nin15_4 nin15 1m
XDIFFw16_p4 sp16_p4 sn16_p4 nin16_4 diff2
Rconn16_p4 nin16_4 nin16 1m
XDIFFw17_p4 sp17_p4 sn17_p4 nin17_4 diff2
Rconn17_p4 nin17_4 nin17 1m
XDIFFw18_p4 sp18_p4 sn18_p4 nin18_4 diff2
Rconn18_p4 nin18_4 nin18 1m
XDIFFw19_p4 sp19_p4 sn19_p4 nin19_4 diff2
Rconn19_p4 nin19_4 nin19 1m
XDIFFw20_p4 sp20_p4 sn20_p4 nin20_4 diff2
Rconn20_p4 nin20_4 nin20 1m
XDIFFw21_p4 sp21_p4 sn21_p4 nin21_4 diff2
Rconn21_p4 nin21_4 nin21 1m
XDIFFw22_p4 sp22_p4 sn22_p4 nin22_4 diff2
Rconn22_p4 nin22_4 nin22 1m
XDIFFw23_p4 sp23_p4 sn23_p4 nin23_4 diff2
Rconn23_p4 nin23_4 nin23 1m
XDIFFw24_p4 sp24_p4 sn24_p4 nin24_4 diff2
Rconn24_p4 nin24_4 nin24 1m
XDIFFw25_p4 sp25_p4 sn25_p4 nin25_4 diff2
Rconn25_p4 nin25_4 nin25 1m
XDIFFw26_p4 sp26_p4 sn26_p4 nin26_4 diff2
Rconn26_p4 nin26_4 nin26 1m
XDIFFw27_p4 sp27_p4 sn27_p4 nin27_4 diff2
Rconn27_p4 nin27_4 nin27 1m
XDIFFw28_p4 sp28_p4 sn28_p4 nin28_4 diff2
Rconn28_p4 nin28_4 nin28 1m
XDIFFw29_p4 sp29_p4 sn29_p4 nin29_4 diff2
Rconn29_p4 nin29_4 nin29 1m
XDIFFw30_p4 sp30_p4 sn30_p4 nin30_4 diff2
Rconn30_p4 nin30_4 nin30 1m
XDIFFw31_p4 sp31_p4 sn31_p4 nin31_4 diff2
Rconn31_p4 nin31_4 nin31 1m
XDIFFw32_p4 sp32_p4 sn32_p4 nin32_4 diff2
Rconn32_p4 nin32_4 nin32 1m
XDIFFw33_p4 sp33_p4 sn33_p4 nin33_4 diff2
Rconn33_p4 nin33_4 nin33 1m
XDIFFw34_p4 sp34_p4 sn34_p4 nin34_4 diff2
Rconn34_p4 nin34_4 nin34 1m
XDIFFw35_p4 sp35_p4 sn35_p4 nin35_4 diff2
Rconn35_p4 nin35_4 nin35 1m
XDIFFw36_p4 sp36_p4 sn36_p4 nin36_4 diff2
Rconn36_p4 nin36_4 nin36 1m
XDIFFw37_p4 sp37_p4 sn37_p4 nin37_4 diff2
Rconn37_p4 nin37_4 nin37 1m
XDIFFw38_p4 sp38_p4 sn38_p4 nin38_4 diff2
Rconn38_p4 nin38_4 nin38 1m
XDIFFw39_p4 sp39_p4 sn39_p4 nin39_4 diff2
Rconn39_p4 nin39_4 nin39 1m
XDIFFw40_p4 sp40_p4 sn40_p4 nin40_4 diff2
Rconn40_p4 nin40_4 nin40 1m
XDIFFw41_p4 sp41_p4 sn41_p4 nin41_4 diff2
Rconn41_p4 nin41_4 nin41 1m
XDIFFw42_p4 sp42_p4 sn42_p4 nin42_4 diff2
Rconn42_p4 nin42_4 nin42 1m
XDIFFw43_p4 sp43_p4 sn43_p4 nin43_4 diff2
Rconn43_p4 nin43_4 nin43 1m
XDIFFw44_p4 sp44_p4 sn44_p4 nin44_4 diff2
Rconn44_p4 nin44_4 nin44 1m
XDIFFw45_p4 sp45_p4 sn45_p4 nin45_4 diff2
Rconn45_p4 nin45_4 nin45 1m
XDIFFw46_p4 sp46_p4 sn46_p4 nin46_4 diff2
Rconn46_p4 nin46_4 nin46 1m
XDIFFw47_p4 sp47_p4 sn47_p4 nin47_4 diff2
Rconn47_p4 nin47_4 nin47 1m
XDIFFw48_p4 sp48_p4 sn48_p4 nin48_4 diff2
Rconn48_p4 nin48_4 nin48 1m
XDIFFw49_p4 sp49_p4 sn49_p4 nin49_4 diff2
Rconn49_p4 nin49_4 nin49 1m
XDIFFw50_p4 sp50_p4 sn50_p4 nin50_4 diff2
Rconn50_p4 nin50_4 nin50 1m
XDIFFw51_p4 sp51_p4 sn51_p4 nin51_4 diff2
Rconn51_p4 nin51_4 nin51 1m
XDIFFw52_p4 sp52_p4 sn52_p4 nin52_4 diff2
Rconn52_p4 nin52_4 nin52 1m
XDIFFw53_p4 sp53_p4 sn53_p4 nin53_4 diff2
Rconn53_p4 nin53_4 nin53 1m
XDIFFw54_p4 sp54_p4 sn54_p4 nin54_4 diff2
Rconn54_p4 nin54_4 nin54 1m
XDIFFw55_p4 sp55_p4 sn55_p4 nin55_4 diff2
Rconn55_p4 nin55_4 nin55 1m
XDIFFw56_p4 sp56_p4 sn56_p4 nin56_4 diff2
Rconn56_p4 nin56_4 nin56 1m
XDIFFw57_p4 sp57_p4 sn57_p4 nin57_4 diff2
Rconn57_p4 nin57_4 nin57 1m
XDIFFw58_p4 sp58_p4 sn58_p4 nin58_4 diff2
Rconn58_p4 nin58_4 nin58 1m
XDIFFw59_p4 sp59_p4 sn59_p4 nin59_4 diff2
Rconn59_p4 nin59_4 nin59 1m
XDIFFw60_p4 sp60_p4 sn60_p4 nin60_4 diff2
Rconn60_p4 nin60_4 nin60 1m
XDIFFw61_p4 sp61_p4 sn61_p4 nin61_4 diff2
Rconn61_p4 nin61_4 nin61 1m
XDIFFw62_p4 sp62_p4 sn62_p4 nin62_4 diff2
Rconn62_p4 nin62_4 nin62 1m
XDIFFw63_p4 sp63_p4 sn63_p4 nin63_4 diff2
Rconn63_p4 nin63_4 nin63 1m
XDIFFw64_p4 sp64_p4 sn64_p4 nin64_4 diff2
Rconn64_p4 nin64_4 nin64 1m
XDIFFw65_p4 sp65_p4 sn65_p4 nin65_4 diff2
Rconn65_p4 nin65_4 nin65 1m
XDIFFw66_p4 sp66_p4 sn66_p4 nin66_4 diff2
Rconn66_p4 nin66_4 nin66 1m
XDIFFw67_p4 sp67_p4 sn67_p4 nin67_4 diff2
Rconn67_p4 nin67_4 nin67 1m
XDIFFw68_p4 sp68_p4 sn68_p4 nin68_4 diff2
Rconn68_p4 nin68_4 nin68 1m
XDIFFw69_p4 sp69_p4 sn69_p4 nin69_4 diff2
Rconn69_p4 nin69_4 nin69 1m
XDIFFw70_p4 sp70_p4 sn70_p4 nin70_4 diff2
Rconn70_p4 nin70_4 nin70 1m
XDIFFw71_p4 sp71_p4 sn71_p4 nin71_4 diff2
Rconn71_p4 nin71_4 nin71 1m
XDIFFw72_p4 sp72_p4 sn72_p4 nin72_4 diff2
Rconn72_p4 nin72_4 nin72 1m
XDIFFw73_p4 sp73_p4 sn73_p4 nin73_4 diff2
Rconn73_p4 nin73_4 nin73 1m
XDIFFw74_p4 sp74_p4 sn74_p4 nin74_4 diff2
Rconn74_p4 nin74_4 nin74 1m
XDIFFw75_p4 sp75_p4 sn75_p4 nin75_4 diff2
Rconn75_p4 nin75_4 nin75 1m
XDIFFw76_p4 sp76_p4 sn76_p4 nin76_4 diff2
Rconn76_p4 nin76_4 nin76 1m
XDIFFw77_p4 sp77_p4 sn77_p4 nin77_4 diff2
Rconn77_p4 nin77_4 nin77 1m
XDIFFw78_p4 sp78_p4 sn78_p4 nin78_4 diff2
Rconn78_p4 nin78_4 nin78 1m
XDIFFw79_p4 sp79_p4 sn79_p4 nin79_4 diff2
Rconn79_p4 nin79_4 nin79 1m
XDIFFw80_p4 sp80_p4 sn80_p4 nin80_4 diff2
Rconn80_p4 nin80_4 nin80 1m
XDIFFw81_p4 sp81_p4 sn81_p4 nin81_4 diff2
Rconn81_p4 nin81_4 nin81 1m
XDIFFw82_p4 sp82_p4 sn82_p4 nin82_4 diff2
Rconn82_p4 nin82_4 nin82 1m
XDIFFw83_p4 sp83_p4 sn83_p4 nin83_4 diff2
Rconn83_p4 nin83_4 nin83 1m
XDIFFw84_p4 sp84_p4 sn84_p4 nin84_4 diff2
Rconn84_p4 nin84_4 nin84 1m


**********neurons****************

Xsig1 nin1 out1 vdd 0 neuron
Xsig2 nin2 out2 vdd 0 neuron
Xsig3 nin3 out3 vdd 0 neuron
Xsig4 nin4 out4 vdd 0 neuron
Xsig5 nin5 out5 vdd 0 neuron
Xsig6 nin6 out6 vdd 0 neuron
Xsig7 nin7 out7 vdd 0 neuron
Xsig8 nin8 out8 vdd 0 neuron
Xsig9 nin9 out9 vdd 0 neuron
Xsig10 nin10 out10 vdd 0 neuron
Xsig11 nin11 out11 vdd 0 neuron
Xsig12 nin12 out12 vdd 0 neuron
Xsig13 nin13 out13 vdd 0 neuron
Xsig14 nin14 out14 vdd 0 neuron
Xsig15 nin15 out15 vdd 0 neuron
Xsig16 nin16 out16 vdd 0 neuron
Xsig17 nin17 out17 vdd 0 neuron
Xsig18 nin18 out18 vdd 0 neuron
Xsig19 nin19 out19 vdd 0 neuron
Xsig20 nin20 out20 vdd 0 neuron
Xsig21 nin21 out21 vdd 0 neuron
Xsig22 nin22 out22 vdd 0 neuron
Xsig23 nin23 out23 vdd 0 neuron
Xsig24 nin24 out24 vdd 0 neuron
Xsig25 nin25 out25 vdd 0 neuron
Xsig26 nin26 out26 vdd 0 neuron
Xsig27 nin27 out27 vdd 0 neuron
Xsig28 nin28 out28 vdd 0 neuron
Xsig29 nin29 out29 vdd 0 neuron
Xsig30 nin30 out30 vdd 0 neuron
Xsig31 nin31 out31 vdd 0 neuron
Xsig32 nin32 out32 vdd 0 neuron
Xsig33 nin33 out33 vdd 0 neuron
Xsig34 nin34 out34 vdd 0 neuron
Xsig35 nin35 out35 vdd 0 neuron
Xsig36 nin36 out36 vdd 0 neuron
Xsig37 nin37 out37 vdd 0 neuron
Xsig38 nin38 out38 vdd 0 neuron
Xsig39 nin39 out39 vdd 0 neuron
Xsig40 nin40 out40 vdd 0 neuron
Xsig41 nin41 out41 vdd 0 neuron
Xsig42 nin42 out42 vdd 0 neuron
Xsig43 nin43 out43 vdd 0 neuron
Xsig44 nin44 out44 vdd 0 neuron
Xsig45 nin45 out45 vdd 0 neuron
Xsig46 nin46 out46 vdd 0 neuron
Xsig47 nin47 out47 vdd 0 neuron
Xsig48 nin48 out48 vdd 0 neuron
Xsig49 nin49 out49 vdd 0 neuron
Xsig50 nin50 out50 vdd 0 neuron
Xsig51 nin51 out51 vdd 0 neuron
Xsig52 nin52 out52 vdd 0 neuron
Xsig53 nin53 out53 vdd 0 neuron
Xsig54 nin54 out54 vdd 0 neuron
Xsig55 nin55 out55 vdd 0 neuron
Xsig56 nin56 out56 vdd 0 neuron
Xsig57 nin57 out57 vdd 0 neuron
Xsig58 nin58 out58 vdd 0 neuron
Xsig59 nin59 out59 vdd 0 neuron
Xsig60 nin60 out60 vdd 0 neuron
Xsig61 nin61 out61 vdd 0 neuron
Xsig62 nin62 out62 vdd 0 neuron
Xsig63 nin63 out63 vdd 0 neuron
Xsig64 nin64 out64 vdd 0 neuron
Xsig65 nin65 out65 vdd 0 neuron
Xsig66 nin66 out66 vdd 0 neuron
Xsig67 nin67 out67 vdd 0 neuron
Xsig68 nin68 out68 vdd 0 neuron
Xsig69 nin69 out69 vdd 0 neuron
Xsig70 nin70 out70 vdd 0 neuron
Xsig71 nin71 out71 vdd 0 neuron
Xsig72 nin72 out72 vdd 0 neuron
Xsig73 nin73 out73 vdd 0 neuron
Xsig74 nin74 out74 vdd 0 neuron
Xsig75 nin75 out75 vdd 0 neuron
Xsig76 nin76 out76 vdd 0 neuron
Xsig77 nin77 out77 vdd 0 neuron
Xsig78 nin78 out78 vdd 0 neuron
Xsig79 nin79 out79 vdd 0 neuron
Xsig80 nin80 out80 vdd 0 neuron
Xsig81 nin81 out81 vdd 0 neuron
Xsig82 nin82 out82 vdd 0 neuron
Xsig83 nin83 out83 vdd 0 neuron
Xsig84 nin84 out84 vdd 0 neuron
.ENDS layer2